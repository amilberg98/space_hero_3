library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity background is
  port(
			clk     : in std_logic;
			y       : in std_logic_vector(9 downto 2);
			x       : in std_logic_vector(9 downto 2);
    		rgb     : out std_logic_vector(5 downto 0)
  	 );
end background;

architecture synth of background is 

	signal address : std_logic_vector(15 downto 0);

begin

		address <= y & x;

		process(clk) begin
			if rising_edge(clk) then
			  case address is
                    when "0000000000110111" => rgb <= "010100";
                    when "0000010001100101" => rgb <= "010100";
                    when "0000010010001100" => rgb <= "000100";
                    when "0000010010001101" => rgb <= "000100";
                    when "0000010101010000" => rgb <= "010100";
                    when "0000011001010000" => rgb <= "010100";
                    when "0001000000000001" => rgb <= "010000";
                    when "0001001001011101" => rgb <= "000100";
                    when "0001001100011100" => rgb <= "010000";
                    when "0001001101011011" => rgb <= "010100";
                    when "0001001101011100" => rgb <= "010100";
                    when "0001001101011101" => rgb <= "000100";
                    when "0001010001011011" => rgb <= "000100";
                    when "0001010001011100" => rgb <= "010100";
                    when "0001010100011011" => rgb <= "010000";
                    when "0001011000100111" => rgb <= "010101";
                    when "0001011001110000" => rgb <= "010000";
                    when "0001011110000110" => rgb <= "010000";
                    when "0001100010000110" => rgb <= "100001";
                    when "0001100010000111" => rgb <= "010000";
                    when "0001110010001000" => rgb <= "010000";
                    when "0001110101011001" => rgb <= "010101";
                    when "0001111000010001" => rgb <= "010000";
                    when "0001111101101110" => rgb <= "101010";
                    when "0001111101101111" => rgb <= "111111";
                    when "0010000001101001" => rgb <= "010101";
                    when "0010100001010101" => rgb <= "010100";
                    when "0010100001010110" => rgb <= "000100";
                    when "0010101001100110" => rgb <= "010000";
                    when "0010101010001100" => rgb <= "010100";
                    when "0010101010001101" => rgb <= "010100";
                    when "0010101010001110" => rgb <= "010100";
                    when "0010101101000100" => rgb <= "000100";
                    when "0010101101000110" => rgb <= "000100";
                    when "0010101101000111" => rgb <= "010100";
                    when "0010101110001100" => rgb <= "010100";
                    when "0010101110001101" => rgb <= "010100";
                    when "0010101110001110" => rgb <= "010100";
                    when "0010110001000111" => rgb <= "000100";
                    when "0010110010001101" => rgb <= "000100";
                    when "0010110100001101" => rgb <= "010000";
                    when "0010111101010101" => rgb <= "000100";
                    when "0010111101101101" => rgb <= "000100";
                    when "0010111110001111" => rgb <= "000100";
                    when "0011000110001001" => rgb <= "011000";
                    when "0011001001101100" => rgb <= "000010";
                    when "0011001101010101" => rgb <= "000100";
                    when "0011001110000010" => rgb <= "000001";
                    when "0011011001111100" => rgb <= "010101";
                    when "0011011010001001" => rgb <= "010000";
                    when "0011011100000110" => rgb <= "011000";
                    when "0011011100000111" => rgb <= "011000";
                    when "0011011100001000" => rgb <= "011000";
                    when "0011100000000110" => rgb <= "011000";
                    when "0011100000000111" => rgb <= "011000";
                    when "0011100000001000" => rgb <= "011000";
                    when "0011100100000111" => rgb <= "010100";
                    when "0011100110001111" => rgb <= "000100";
                    when "0011100110010000" => rgb <= "000100";
                    when "0011101000110000" => rgb <= "100001";
                    when "0011101000110110" => rgb <= "010000";
                    when "0011101010001110" => rgb <= "000100";
                    when "0011101010010000" => rgb <= "000100";
                    when "0011101010010010" => rgb <= "011000";
                    when "0011101100100101" => rgb <= "010000";
                    when "0011101101011011" => rgb <= "000100";
                    when "0011101110010000" => rgb <= "000100";
                    when "0011101110010010" => rgb <= "011000";
                    when "0011101110010011" => rgb <= "010100";
                    when "0011110000100010" => rgb <= "010101";
                    when "0011110010010000" => rgb <= "000100";
                    when "0011110010010010" => rgb <= "011000";
                    when "0011110110010010" => rgb <= "000100";
                    when "0011111001101110" => rgb <= "000100";
                    when "0011111001101111" => rgb <= "010100";
                    when "0011111001110000" => rgb <= "010101";
                    when "0011111101101110" => rgb <= "010100";
                    when "0011111101101111" => rgb <= "010101";
                    when "0011111101110000" => rgb <= "011000";
                    when "0011111101110001" => rgb <= "010100";
                    when "0100000001101110" => rgb <= "010100";
                    when "0100000001101111" => rgb <= "011000";
                    when "0100000001110000" => rgb <= "011000";
                    when "0100000001110001" => rgb <= "010100";
                    when "0100000001110011" => rgb <= "000110";
                    when "0100000101101111" => rgb <= "010100";
                    when "0100000101110000" => rgb <= "010100";
                    when "0100000101110001" => rgb <= "000100";
                    when "0100001000000100" => rgb <= "010000";
                    when "0100001001111100" => rgb <= "010000";
                    when "0100001001111101" => rgb <= "100001";
                    when "0100001001111110" => rgb <= "100001";
                    when "0100001010000110" => rgb <= "000100";
                    when "0100001101111100" => rgb <= "100001";
                    when "0100001101111101" => rgb <= "100001";
                    when "0100001101111110" => rgb <= "100001";
                    when "0100001110000110" => rgb <= "000100";
                    when "0100010000100111" => rgb <= "101010";
                    when "0100010000101000" => rgb <= "101010";
                    when "0100011101100010" => rgb <= "000100";
                    when "0100100000000110" => rgb <= "010100";
                    when "0100101000001110" => rgb <= "010000";
                    when "0100110001000100" => rgb <= "011000";
                    when "0100110001000101" => rgb <= "000100";
                    when "0100110100101111" => rgb <= "010000";
                    when "0100110101000100" => rgb <= "011000";
                    when "0100110101000101" => rgb <= "010100";
                    when "0100111110000101" => rgb <= "010100";
                    when "0100111110001000" => rgb <= "010100";
                    when "0100111110001001" => rgb <= "010100";
                    when "0100111110001010" => rgb <= "010100";
                    when "0101000010001000" => rgb <= "010100";
                    when "0101000010001001" => rgb <= "010100";
                    when "0101000100101001" => rgb <= "000001";
                    when "0101000100101010" => rgb <= "000010";
                    when "0101010100110011" => rgb <= "000100";
                    when "0101010110000000" => rgb <= "010100";
                    when "0101010110000001" => rgb <= "011000";
                    when "0101010110000011" => rgb <= "010100";
                    when "0101011000110011" => rgb <= "000100";
                    when "0101011010011110" => rgb <= "010100";
                    when "0101011010011111" => rgb <= "010100";
                    when "0101011101000010" => rgb <= "010100";
                    when "0101011101000011" => rgb <= "010100";
                    when "0101011110011111" => rgb <= "010100";
                    when "0101100001000010" => rgb <= "000100";
                    when "0101100001000011" => rgb <= "010100";
                    when "0101101000100100" => rgb <= "010000";
                    when "0101101100110111" => rgb <= "010100";
                    when "0101101100111000" => rgb <= "010100";
                    when "0101101101001000" => rgb <= "010100";
                    when "0101110001000110" => rgb <= "000100";
                    when "0101111000001101" => rgb <= "010100";
                    when "0101111000001110" => rgb <= "000100";
                    when "0101111001111010" => rgb <= "000100";
                    when "0101111001111011" => rgb <= "000100";
                    when "0101111100001110" => rgb <= "000100";
                    when "0110000000001100" => rgb <= "000100";
                    when "0110000000001110" => rgb <= "000100";
                    when "0110000101011011" => rgb <= "000100";
                    when "0110000101011100" => rgb <= "010100";
                    when "0110000101011101" => rgb <= "010100";
                    when "0110001001011011" => rgb <= "010100";
                    when "0110001001011100" => rgb <= "010100";
                    when "0110001001011101" => rgb <= "010100";
                    when "0110001001011110" => rgb <= "000100";
                    when "0110001100000000" => rgb <= "101010";
                    when "0110001100000001" => rgb <= "101010";
                    when "0110001100000100" => rgb <= "101010";
                    when "0110001100001010" => rgb <= "101010";
                    when "0110001100001110" => rgb <= "101010";
                    when "0110001100010000" => rgb <= "101010";
                    when "0110001100010001" => rgb <= "101010";
                    when "0110001100010111" => rgb <= "101010";
                    when "0110001100100000" => rgb <= "101010";
                    when "0110001100100001" => rgb <= "101010";
                    when "0110001100100110" => rgb <= "101010";
                    when "0110001100101001" => rgb <= "101010";
                    when "0110001100110000" => rgb <= "101010";
                    when "0110001100110001" => rgb <= "101010";
                    when "0110001100111101" => rgb <= "101010";
                    when "0110001101000000" => rgb <= "101010";
                    when "0110001101000001" => rgb <= "101010";
                    when "0110001101000100" => rgb <= "101010";
                    when "0110001101001010" => rgb <= "101010";
                    when "0110001101001011" => rgb <= "010100";
                    when "0110001101001100" => rgb <= "010100";
                    when "0110001101001101" => rgb <= "010100";
                    when "0110001101001110" => rgb <= "101010";
                    when "0110001101001111" => rgb <= "010100";
                    when "0110001101010000" => rgb <= "101010";
                    when "0110001101010001" => rgb <= "101010";
                    when "0110001101010111" => rgb <= "101010";
                    when "0110001101011011" => rgb <= "000100";
                    when "0110001101011100" => rgb <= "010100";
                    when "0110001101011101" => rgb <= "010100";
                    when "0110001101100000" => rgb <= "101010";
                    when "0110001101100001" => rgb <= "101010";
                    when "0110001101100110" => rgb <= "101010";
                    when "0110001101101001" => rgb <= "101010";
                    when "0110001101110000" => rgb <= "101010";
                    when "0110001101110001" => rgb <= "101010";
                    when "0110001101111101" => rgb <= "101010";
                    when "0110001101111111" => rgb <= "000100";
                    when "0110001110000000" => rgb <= "101010";
                    when "0110001110000001" => rgb <= "101010";
                    when "0110001110000110" => rgb <= "101010";
                    when "0110001110001001" => rgb <= "101010";
                    when "0110001110010000" => rgb <= "101010";
                    when "0110001110010001" => rgb <= "101010";
                    when "0110001110011101" => rgb <= "101010";
                    when "0110010000000000" => rgb <= "101010";
                    when "0110010000000001" => rgb <= "101010";
                    when "0110010000000010" => rgb <= "101010";
                    when "0110010000000011" => rgb <= "101010";
                    when "0110010000000100" => rgb <= "101010";
                    when "0110010000000101" => rgb <= "101010";
                    when "0110010000000110" => rgb <= "101010";
                    when "0110010000000111" => rgb <= "101010";
                    when "0110010000001000" => rgb <= "101010";
                    when "0110010000001001" => rgb <= "101010";
                    when "0110010000001010" => rgb <= "101010";
                    when "0110010000001011" => rgb <= "101010";
                    when "0110010000001100" => rgb <= "101010";
                    when "0110010000001101" => rgb <= "101010";
                    when "0110010000001110" => rgb <= "101010";
                    when "0110010000001111" => rgb <= "101010";
                    when "0110010000010000" => rgb <= "101010";
                    when "0110010000010001" => rgb <= "101010";
                    when "0110010000010010" => rgb <= "101010";
                    when "0110010000010011" => rgb <= "101010";
                    when "0110010000010100" => rgb <= "101010";
                    when "0110010000010101" => rgb <= "101010";
                    when "0110010000010110" => rgb <= "101010";
                    when "0110010000010111" => rgb <= "101010";
                    when "0110010000011000" => rgb <= "101010";
                    when "0110010000011001" => rgb <= "101010";
                    when "0110010000011010" => rgb <= "101010";
                    when "0110010000011011" => rgb <= "101010";
                    when "0110010000011100" => rgb <= "101010";
                    when "0110010000011101" => rgb <= "101010";
                    when "0110010000011110" => rgb <= "101010";
                    when "0110010000011111" => rgb <= "101010";
                    when "0110010000100000" => rgb <= "101010";
                    when "0110010000100001" => rgb <= "101010";
                    when "0110010000100010" => rgb <= "101010";
                    when "0110010000100011" => rgb <= "101010";
                    when "0110010000100100" => rgb <= "101010";
                    when "0110010000100101" => rgb <= "101010";
                    when "0110010000100110" => rgb <= "101010";
                    when "0110010000100111" => rgb <= "101010";
                    when "0110010000101000" => rgb <= "101010";
                    when "0110010000101001" => rgb <= "101010";
                    when "0110010000101010" => rgb <= "101010";
                    when "0110010000101011" => rgb <= "101010";
                    when "0110010000101100" => rgb <= "101010";
                    when "0110010000101101" => rgb <= "101010";
                    when "0110010000101110" => rgb <= "101010";
                    when "0110010000101111" => rgb <= "101010";
                    when "0110010000110000" => rgb <= "101010";
                    when "0110010000110001" => rgb <= "101010";
                    when "0110010000110010" => rgb <= "101010";
                    when "0110010000110011" => rgb <= "101010";
                    when "0110010000110100" => rgb <= "101010";
                    when "0110010000110101" => rgb <= "101010";
                    when "0110010000110110" => rgb <= "101010";
                    when "0110010000110111" => rgb <= "101010";
                    when "0110010000111000" => rgb <= "101010";
                    when "0110010000111001" => rgb <= "101010";
                    when "0110010000111010" => rgb <= "101010";
                    when "0110010000111011" => rgb <= "101010";
                    when "0110010000111100" => rgb <= "101010";
                    when "0110010000111101" => rgb <= "101010";
                    when "0110010000111110" => rgb <= "101010";
                    when "0110010000111111" => rgb <= "101010";
                    when "0110010001000000" => rgb <= "101010";
                    when "0110010001000001" => rgb <= "101010";
                    when "0110010001000010" => rgb <= "101010";
                    when "0110010001000011" => rgb <= "101010";
                    when "0110010001000100" => rgb <= "101010";
                    when "0110010001000101" => rgb <= "101010";
                    when "0110010001000110" => rgb <= "101010";
                    when "0110010001000111" => rgb <= "101010";
                    when "0110010001001000" => rgb <= "101010";
                    when "0110010001001001" => rgb <= "101010";
                    when "0110010001001010" => rgb <= "101010";
                    when "0110010001001011" => rgb <= "101010";
                    when "0110010001001100" => rgb <= "101010";
                    when "0110010001001101" => rgb <= "101010";
                    when "0110010001001110" => rgb <= "101010";
                    when "0110010001001111" => rgb <= "101010";
                    when "0110010001010000" => rgb <= "101010";
                    when "0110010001010001" => rgb <= "101010";
                    when "0110010001010010" => rgb <= "101010";
                    when "0110010001010011" => rgb <= "101010";
                    when "0110010001010100" => rgb <= "101010";
                    when "0110010001010101" => rgb <= "101010";
                    when "0110010001010110" => rgb <= "101010";
                    when "0110010001010111" => rgb <= "101010";
                    when "0110010001011000" => rgb <= "101010";
                    when "0110010001011001" => rgb <= "101010";
                    when "0110010001011010" => rgb <= "101010";
                    when "0110010001011011" => rgb <= "101010";
                    when "0110010001011100" => rgb <= "101010";
                    when "0110010001011101" => rgb <= "101010";
                    when "0110010001011110" => rgb <= "101010";
                    when "0110010001011111" => rgb <= "101010";
                    when "0110010001100000" => rgb <= "101010";
                    when "0110010001100001" => rgb <= "101010";
                    when "0110010001100010" => rgb <= "101010";
                    when "0110010001100011" => rgb <= "101010";
                    when "0110010001100100" => rgb <= "101010";
                    when "0110010001100101" => rgb <= "101010";
                    when "0110010001100110" => rgb <= "101010";
                    when "0110010001100111" => rgb <= "101010";
                    when "0110010001101000" => rgb <= "101010";
                    when "0110010001101001" => rgb <= "101010";
                    when "0110010001101010" => rgb <= "101010";
                    when "0110010001101011" => rgb <= "101010";
                    when "0110010001101100" => rgb <= "101010";
                    when "0110010001101101" => rgb <= "101010";
                    when "0110010001101110" => rgb <= "101010";
                    when "0110010001101111" => rgb <= "101010";
                    when "0110010001110000" => rgb <= "101010";
                    when "0110010001110001" => rgb <= "101010";
                    when "0110010001110010" => rgb <= "101010";
                    when "0110010001110011" => rgb <= "101010";
                    when "0110010001110100" => rgb <= "101010";
                    when "0110010001110101" => rgb <= "101010";
                    when "0110010001110110" => rgb <= "101010";
                    when "0110010001110111" => rgb <= "101010";
                    when "0110010001111000" => rgb <= "101010";
                    when "0110010001111001" => rgb <= "101010";
                    when "0110010001111010" => rgb <= "101010";
                    when "0110010001111011" => rgb <= "101010";
                    when "0110010001111100" => rgb <= "101010";
                    when "0110010001111101" => rgb <= "101010";
                    when "0110010001111110" => rgb <= "101010";
                    when "0110010001111111" => rgb <= "101010";
                    when "0110010010000000" => rgb <= "101010";
                    when "0110010010000001" => rgb <= "101010";
                    when "0110010010000010" => rgb <= "101010";
                    when "0110010010000011" => rgb <= "101010";
                    when "0110010010000100" => rgb <= "101010";
                    when "0110010010000101" => rgb <= "101010";
                    when "0110010010000110" => rgb <= "101010";
                    when "0110010010000111" => rgb <= "101010";
                    when "0110010010001000" => rgb <= "101010";
                    when "0110010010001001" => rgb <= "101010";
                    when "0110010010001010" => rgb <= "101010";
                    when "0110010010001011" => rgb <= "101010";
                    when "0110010010001100" => rgb <= "101010";
                    when "0110010010001101" => rgb <= "101010";
                    when "0110010010001110" => rgb <= "101010";
                    when "0110010010001111" => rgb <= "101010";
                    when "0110010010010000" => rgb <= "101010";
                    when "0110010010010001" => rgb <= "101010";
                    when "0110010010010010" => rgb <= "101010";
                    when "0110010010010011" => rgb <= "101010";
                    when "0110010010010100" => rgb <= "101010";
                    when "0110010010010101" => rgb <= "101010";
                    when "0110010010010110" => rgb <= "101010";
                    when "0110010010010111" => rgb <= "101010";
                    when "0110010010011000" => rgb <= "101010";
                    when "0110010010011001" => rgb <= "101010";
                    when "0110010010011010" => rgb <= "101010";
                    when "0110010010011011" => rgb <= "101010";
                    when "0110010010011100" => rgb <= "101010";
                    when "0110010010011101" => rgb <= "101010";
                    when "0110010010011110" => rgb <= "101010";
                    when "0110010010011111" => rgb <= "101010";
                    when "0110010100000000" => rgb <= "101010";
                    when "0110010100000001" => rgb <= "101010";
                    when "0110010100010000" => rgb <= "101010";
                    when "0110010100010001" => rgb <= "101010";
                    when "0110010100100000" => rgb <= "101010";
                    when "0110010100100001" => rgb <= "101010";
                    when "0110010100110000" => rgb <= "101010";
                    when "0110010100110001" => rgb <= "101010";
                    when "0110010101000000" => rgb <= "101010";
                    when "0110010101000001" => rgb <= "101010";
                    when "0110010101010000" => rgb <= "101010";
                    when "0110010101010001" => rgb <= "101010";
                    when "0110010101100000" => rgb <= "101010";
                    when "0110010101100001" => rgb <= "101010";
                    when "0110010101110000" => rgb <= "101010";
                    when "0110010101110001" => rgb <= "101010";
                    when "0110010110000000" => rgb <= "101010";
                    when "0110010110000001" => rgb <= "101010";
                    when "0110010110010000" => rgb <= "101010";
                    when "0110010110010001" => rgb <= "101010";
                    when "0110011000000000" => rgb <= "010101";
                    when "0110011000000001" => rgb <= "010101";
                    when "0110011000000010" => rgb <= "010101";
                    when "0110011000000011" => rgb <= "010101";
                    when "0110011000000100" => rgb <= "010101";
                    when "0110011000000101" => rgb <= "010101";
                    when "0110011000000110" => rgb <= "010101";
                    when "0110011000000111" => rgb <= "010101";
                    when "0110011000001000" => rgb <= "010101";
                    when "0110011000001001" => rgb <= "010101";
                    when "0110011000001010" => rgb <= "010101";
                    when "0110011000001011" => rgb <= "010101";
                    when "0110011000001100" => rgb <= "010101";
                    when "0110011000001101" => rgb <= "010101";
                    when "0110011000001110" => rgb <= "010101";
                    when "0110011000001111" => rgb <= "010101";
                    when "0110011000010000" => rgb <= "010101";
                    when "0110011000010001" => rgb <= "010101";
                    when "0110011000010010" => rgb <= "010101";
                    when "0110011000010011" => rgb <= "010101";
                    when "0110011000010100" => rgb <= "010101";
                    when "0110011000010101" => rgb <= "010101";
                    when "0110011000010110" => rgb <= "010101";
                    when "0110011000010111" => rgb <= "010101";
                    when "0110011000011000" => rgb <= "010101";
                    when "0110011000011001" => rgb <= "010101";
                    when "0110011000011010" => rgb <= "010101";
                    when "0110011000011011" => rgb <= "010101";
                    when "0110011000011100" => rgb <= "010101";
                    when "0110011000011101" => rgb <= "010101";
                    when "0110011000011110" => rgb <= "010101";
                    when "0110011000011111" => rgb <= "010101";
                    when "0110011000100000" => rgb <= "010101";
                    when "0110011000100001" => rgb <= "010101";
                    when "0110011000100010" => rgb <= "010101";
                    when "0110011000100011" => rgb <= "010101";
                    when "0110011000100100" => rgb <= "010101";
                    when "0110011000100101" => rgb <= "010101";
                    when "0110011000100110" => rgb <= "010101";
                    when "0110011000100111" => rgb <= "010101";
                    when "0110011000101000" => rgb <= "010101";
                    when "0110011000101001" => rgb <= "010101";
                    when "0110011000101010" => rgb <= "010101";
                    when "0110011000101011" => rgb <= "010101";
                    when "0110011000101100" => rgb <= "010101";
                    when "0110011000101101" => rgb <= "010101";
                    when "0110011000101110" => rgb <= "010101";
                    when "0110011000101111" => rgb <= "010101";
                    when "0110011000110000" => rgb <= "010101";
                    when "0110011000110001" => rgb <= "010101";
                    when "0110011000110010" => rgb <= "010101";
                    when "0110011000110011" => rgb <= "010101";
                    when "0110011000110100" => rgb <= "010101";
                    when "0110011000110101" => rgb <= "010101";
                    when "0110011000110110" => rgb <= "010101";
                    when "0110011000110111" => rgb <= "010101";
                    when "0110011000111000" => rgb <= "010101";
                    when "0110011000111001" => rgb <= "010101";
                    when "0110011000111010" => rgb <= "010101";
                    when "0110011000111011" => rgb <= "010101";
                    when "0110011000111100" => rgb <= "010101";
                    when "0110011000111101" => rgb <= "010101";
                    when "0110011000111110" => rgb <= "010101";
                    when "0110011000111111" => rgb <= "010101";
                    when "0110011001000000" => rgb <= "010101";
                    when "0110011001000001" => rgb <= "010101";
                    when "0110011001000010" => rgb <= "010101";
                    when "0110011001000011" => rgb <= "010101";
                    when "0110011001000100" => rgb <= "010101";
                    when "0110011001000101" => rgb <= "010101";
                    when "0110011001000110" => rgb <= "010101";
                    when "0110011001000111" => rgb <= "010101";
                    when "0110011001001000" => rgb <= "010101";
                    when "0110011001001001" => rgb <= "010101";
                    when "0110011001001010" => rgb <= "010101";
                    when "0110011001001011" => rgb <= "010101";
                    when "0110011001001100" => rgb <= "010101";
                    when "0110011001001101" => rgb <= "010101";
                    when "0110011001001110" => rgb <= "010101";
                    when "0110011001001111" => rgb <= "010101";
                    when "0110011001010000" => rgb <= "010101";
                    when "0110011001010001" => rgb <= "010101";
                    when "0110011001010010" => rgb <= "010101";
                    when "0110011001010011" => rgb <= "010101";
                    when "0110011001010100" => rgb <= "010101";
                    when "0110011001010101" => rgb <= "010101";
                    when "0110011001010110" => rgb <= "010101";
                    when "0110011001010111" => rgb <= "010101";
                    when "0110011001011000" => rgb <= "010101";
                    when "0110011001011001" => rgb <= "010101";
                    when "0110011001011010" => rgb <= "010101";
                    when "0110011001011011" => rgb <= "010101";
                    when "0110011001011100" => rgb <= "010101";
                    when "0110011001011101" => rgb <= "010101";
                    when "0110011001011110" => rgb <= "010101";
                    when "0110011001011111" => rgb <= "010101";
                    when "0110011001100000" => rgb <= "010101";
                    when "0110011001100001" => rgb <= "010101";
                    when "0110011001100010" => rgb <= "010101";
                    when "0110011001100011" => rgb <= "010101";
                    when "0110011001100100" => rgb <= "010101";
                    when "0110011001100101" => rgb <= "010101";
                    when "0110011001100110" => rgb <= "010101";
                    when "0110011001100111" => rgb <= "010101";
                    when "0110011001101000" => rgb <= "010101";
                    when "0110011001101001" => rgb <= "010101";
                    when "0110011001101010" => rgb <= "010101";
                    when "0110011001101011" => rgb <= "010101";
                    when "0110011001101100" => rgb <= "010101";
                    when "0110011001101101" => rgb <= "010101";
                    when "0110011001101110" => rgb <= "010101";
                    when "0110011001101111" => rgb <= "010101";
                    when "0110011001110000" => rgb <= "010101";
                    when "0110011001110001" => rgb <= "010101";
                    when "0110011001110010" => rgb <= "010101";
                    when "0110011001110011" => rgb <= "010101";
                    when "0110011001110100" => rgb <= "010101";
                    when "0110011001110101" => rgb <= "010101";
                    when "0110011001110110" => rgb <= "010101";
                    when "0110011001110111" => rgb <= "010101";
                    when "0110011001111000" => rgb <= "010101";
                    when "0110011001111001" => rgb <= "010101";
                    when "0110011001111010" => rgb <= "010101";
                    when "0110011001111011" => rgb <= "010101";
                    when "0110011001111100" => rgb <= "010101";
                    when "0110011001111101" => rgb <= "010101";
                    when "0110011001111110" => rgb <= "010101";
                    when "0110011001111111" => rgb <= "010101";
                    when "0110011010000000" => rgb <= "010101";
                    when "0110011010000001" => rgb <= "010101";
                    when "0110011010000010" => rgb <= "010101";
                    when "0110011010000011" => rgb <= "010101";
                    when "0110011010000100" => rgb <= "010101";
                    when "0110011010000101" => rgb <= "010101";
                    when "0110011010000110" => rgb <= "010101";
                    when "0110011010000111" => rgb <= "010101";
                    when "0110011010001000" => rgb <= "010101";
                    when "0110011010001001" => rgb <= "010101";
                    when "0110011010001010" => rgb <= "010101";
                    when "0110011010001011" => rgb <= "010101";
                    when "0110011010001100" => rgb <= "010101";
                    when "0110011010001101" => rgb <= "010101";
                    when "0110011010001110" => rgb <= "010101";
                    when "0110011010001111" => rgb <= "010101";
                    when "0110011010010000" => rgb <= "010101";
                    when "0110011010010001" => rgb <= "010101";
                    when "0110011010010010" => rgb <= "010101";
                    when "0110011010010011" => rgb <= "010101";
                    when "0110011010010100" => rgb <= "010101";
                    when "0110011010010101" => rgb <= "010101";
                    when "0110011010010110" => rgb <= "010101";
                    when "0110011010010111" => rgb <= "010101";
                    when "0110011010011000" => rgb <= "010101";
                    when "0110011010011001" => rgb <= "010101";
                    when "0110011010011010" => rgb <= "010101";
                    when "0110011010011011" => rgb <= "010101";
                    when "0110011010011100" => rgb <= "010101";
                    when "0110011010011101" => rgb <= "010101";
                    when "0110011010011110" => rgb <= "010101";
                    when "0110011010011111" => rgb <= "010101";
                    when "0110011100000000" => rgb <= "101010";
                    when "0110011100000001" => rgb <= "101010";
                    when "0110011100010000" => rgb <= "101010";
                    when "0110011100010001" => rgb <= "101010";
                    when "0110011100100000" => rgb <= "101010";
                    when "0110011100100001" => rgb <= "101010";
                    when "0110011100110000" => rgb <= "101010";
                    when "0110011100110001" => rgb <= "101010";
                    when "0110011101000000" => rgb <= "101010";
                    when "0110011101000001" => rgb <= "101010";
                    when "0110011101010000" => rgb <= "101010";
                    when "0110011101010001" => rgb <= "101010";
                    when "0110011101110000" => rgb <= "101010";
                    when "0110011101110001" => rgb <= "101010";
                    when "0110011110000000" => rgb <= "101010";
                    when "0110011110000001" => rgb <= "101010";
                    when "0110011110010000" => rgb <= "101010";
                    when "0110011110010001" => rgb <= "101010";
                    when "0110100000000000" => rgb <= "101010";
                    when "0110100000000001" => rgb <= "101010";
                    when "0110100000000011" => rgb <= "101010";
                    when "0110100000000100" => rgb <= "101010";
                    when "0110100000000101" => rgb <= "101010";
                    when "0110100000000110" => rgb <= "101010";
                    when "0110100000000111" => rgb <= "101010";
                    when "0110100000001000" => rgb <= "101010";
                    when "0110100000001001" => rgb <= "101010";
                    when "0110100000001010" => rgb <= "101010";
                    when "0110100000001011" => rgb <= "101010";
                    when "0110100000001100" => rgb <= "101010";
                    when "0110100000001101" => rgb <= "101010";
                    when "0110100000001110" => rgb <= "101010";
                    when "0110100000010000" => rgb <= "101010";
                    when "0110100000010001" => rgb <= "101010";
                    when "0110100000010011" => rgb <= "101010";
                    when "0110100000010100" => rgb <= "101010";
                    when "0110100000010101" => rgb <= "101010";
                    when "0110100000010110" => rgb <= "101010";
                    when "0110100000010111" => rgb <= "101010";
                    when "0110100000011000" => rgb <= "101010";
                    when "0110100000011001" => rgb <= "101010";
                    when "0110100000011010" => rgb <= "101010";
                    when "0110100000011011" => rgb <= "101010";
                    when "0110100000011100" => rgb <= "101010";
                    when "0110100000011101" => rgb <= "101010";
                    when "0110100000011110" => rgb <= "101010";
                    when "0110100000100000" => rgb <= "101010";
                    when "0110100000100001" => rgb <= "101010";
                    when "0110100000100011" => rgb <= "101010";
                    when "0110100000100100" => rgb <= "101010";
                    when "0110100000100101" => rgb <= "101010";
                    when "0110100000100110" => rgb <= "101010";
                    when "0110100000100111" => rgb <= "101010";
                    when "0110100000101000" => rgb <= "101010";
                    when "0110100000101001" => rgb <= "101010";
                    when "0110100000101010" => rgb <= "101010";
                    when "0110100000101011" => rgb <= "101010";
                    when "0110100000101100" => rgb <= "101010";
                    when "0110100000101101" => rgb <= "101010";
                    when "0110100000101110" => rgb <= "101010";
                    when "0110100000110000" => rgb <= "101010";
                    when "0110100000110001" => rgb <= "101010";
                    when "0110100000110011" => rgb <= "101010";
                    when "0110100000110100" => rgb <= "101010";
                    when "0110100000110101" => rgb <= "101010";
                    when "0110100000110110" => rgb <= "101010";
                    when "0110100000110111" => rgb <= "101010";
                    when "0110100000111000" => rgb <= "101010";
                    when "0110100000111001" => rgb <= "101010";
                    when "0110100000111010" => rgb <= "101010";
                    when "0110100000111011" => rgb <= "101010";
                    when "0110100000111100" => rgb <= "101010";
                    when "0110100000111101" => rgb <= "101010";
                    when "0110100000111110" => rgb <= "101010";
                    when "0110100001000000" => rgb <= "101010";
                    when "0110100001000001" => rgb <= "101010";
                    when "0110100001000011" => rgb <= "101010";
                    when "0110100001000100" => rgb <= "101010";
                    when "0110100001000101" => rgb <= "101010";
                    when "0110100001000110" => rgb <= "101010";
                    when "0110100001000111" => rgb <= "101010";
                    when "0110100001001000" => rgb <= "101010";
                    when "0110100001001001" => rgb <= "101010";
                    when "0110100001001010" => rgb <= "101010";
                    when "0110100001001011" => rgb <= "101010";
                    when "0110100001001100" => rgb <= "101010";
                    when "0110100001001101" => rgb <= "101010";
                    when "0110100001001110" => rgb <= "101010";
                    when "0110100001010000" => rgb <= "101010";
                    when "0110100001010001" => rgb <= "101010";
                    when "0110100001010011" => rgb <= "101010";
                    when "0110100001010100" => rgb <= "101010";
                    when "0110100001010101" => rgb <= "101010";
                    when "0110100001011100" => rgb <= "101010";
                    when "0110100001011101" => rgb <= "101010";
                    when "0110100001011110" => rgb <= "101010";
                    when "0110100001011111" => rgb <= "101010";
                    when "0110100001100000" => rgb <= "101010";
                    when "0110100001100001" => rgb <= "101010";
                    when "0110100001100010" => rgb <= "101010";
                    when "0110100001100011" => rgb <= "101010";
                    when "0110100001100100" => rgb <= "101010";
                    when "0110100001100101" => rgb <= "101010";
                    when "0110100001100110" => rgb <= "101010";
                    when "0110100001100111" => rgb <= "101010";
                    when "0110100001101000" => rgb <= "101010";
                    when "0110100001101001" => rgb <= "101010";
                    when "0110100001101010" => rgb <= "101010";
                    when "0110100001101011" => rgb <= "101010";
                    when "0110100001101100" => rgb <= "101010";
                    when "0110100001101101" => rgb <= "101010";
                    when "0110100001101110" => rgb <= "101010";
                    when "0110100001101111" => rgb <= "101010";
                    when "0110100001110000" => rgb <= "101010";
                    when "0110100001110001" => rgb <= "101010";
                    when "0110100001110011" => rgb <= "101010";
                    when "0110100001110100" => rgb <= "101010";
                    when "0110100001110101" => rgb <= "101010";
                    when "0110100001110110" => rgb <= "101010";
                    when "0110100001110111" => rgb <= "101010";
                    when "0110100001111000" => rgb <= "101010";
                    when "0110100001111001" => rgb <= "101010";
                    when "0110100001111010" => rgb <= "101010";
                    when "0110100001111011" => rgb <= "101010";
                    when "0110100001111100" => rgb <= "101010";
                    when "0110100001111101" => rgb <= "101010";
                    when "0110100001111110" => rgb <= "101010";
                    when "0110100010000000" => rgb <= "101010";
                    when "0110100010000001" => rgb <= "101010";
                    when "0110100010000011" => rgb <= "101010";
                    when "0110100010000100" => rgb <= "101010";
                    when "0110100010000101" => rgb <= "101010";
                    when "0110100010000110" => rgb <= "101010";
                    when "0110100010000111" => rgb <= "101010";
                    when "0110100010001000" => rgb <= "101010";
                    when "0110100010001001" => rgb <= "101010";
                    when "0110100010001010" => rgb <= "101010";
                    when "0110100010001011" => rgb <= "101010";
                    when "0110100010001100" => rgb <= "101010";
                    when "0110100010001101" => rgb <= "101010";
                    when "0110100010001110" => rgb <= "101010";
                    when "0110100010010000" => rgb <= "101010";
                    when "0110100010010001" => rgb <= "101010";
                    when "0110100010010011" => rgb <= "101010";
                    when "0110100010010100" => rgb <= "101010";
                    when "0110100010010101" => rgb <= "101010";
                    when "0110100010010110" => rgb <= "101010";
                    when "0110100010010111" => rgb <= "101010";
                    when "0110100010011000" => rgb <= "101010";
                    when "0110100010011001" => rgb <= "101010";
                    when "0110100010011010" => rgb <= "101010";
                    when "0110100010011011" => rgb <= "101010";
                    when "0110100010011100" => rgb <= "101010";
                    when "0110100010011101" => rgb <= "101010";
                    when "0110100010011110" => rgb <= "101010";
                    when "0110100100000000" => rgb <= "101010";
                    when "0110100100000001" => rgb <= "101010";
                    when "0110100100000011" => rgb <= "010101";
                    when "0110100100000100" => rgb <= "010101";
                    when "0110100100000101" => rgb <= "010101";
                    when "0110100100000110" => rgb <= "010101";
                    when "0110100100000111" => rgb <= "010101";
                    when "0110100100001000" => rgb <= "010101";
                    when "0110100100001001" => rgb <= "010101";
                    when "0110100100001010" => rgb <= "010101";
                    when "0110100100001011" => rgb <= "010101";
                    when "0110100100001100" => rgb <= "010101";
                    when "0110100100001101" => rgb <= "010101";
                    when "0110100100001110" => rgb <= "010101";
                    when "0110100100010000" => rgb <= "101010";
                    when "0110100100010001" => rgb <= "101010";
                    when "0110100100010011" => rgb <= "010101";
                    when "0110100100010100" => rgb <= "010101";
                    when "0110100100010101" => rgb <= "010101";
                    when "0110100100010110" => rgb <= "010101";
                    when "0110100100010111" => rgb <= "010101";
                    when "0110100100011000" => rgb <= "010101";
                    when "0110100100011001" => rgb <= "010101";
                    when "0110100100011010" => rgb <= "010101";
                    when "0110100100011011" => rgb <= "010101";
                    when "0110100100011100" => rgb <= "010101";
                    when "0110100100011101" => rgb <= "010101";
                    when "0110100100011110" => rgb <= "010101";
                    when "0110100100100000" => rgb <= "101010";
                    when "0110100100100001" => rgb <= "101010";
                    when "0110100100100011" => rgb <= "010101";
                    when "0110100100100100" => rgb <= "010101";
                    when "0110100100100101" => rgb <= "010101";
                    when "0110100100100110" => rgb <= "010101";
                    when "0110100100100111" => rgb <= "010101";
                    when "0110100100101000" => rgb <= "010101";
                    when "0110100100101001" => rgb <= "010101";
                    when "0110100100101010" => rgb <= "010101";
                    when "0110100100101011" => rgb <= "010101";
                    when "0110100100101100" => rgb <= "010101";
                    when "0110100100101101" => rgb <= "010101";
                    when "0110100100101110" => rgb <= "010101";
                    when "0110100100110000" => rgb <= "101010";
                    when "0110100100110001" => rgb <= "101010";
                    when "0110100100110011" => rgb <= "010101";
                    when "0110100100110100" => rgb <= "010101";
                    when "0110100100110101" => rgb <= "010101";
                    when "0110100100110110" => rgb <= "010101";
                    when "0110100100110111" => rgb <= "010101";
                    when "0110100100111000" => rgb <= "010101";
                    when "0110100100111001" => rgb <= "010101";
                    when "0110100100111010" => rgb <= "010101";
                    when "0110100100111011" => rgb <= "010101";
                    when "0110100100111100" => rgb <= "010101";
                    when "0110100100111101" => rgb <= "010101";
                    when "0110100100111110" => rgb <= "010101";
                    when "0110100101000000" => rgb <= "101010";
                    when "0110100101000001" => rgb <= "101010";
                    when "0110100101000011" => rgb <= "010101";
                    when "0110100101000100" => rgb <= "010101";
                    when "0110100101000101" => rgb <= "010101";
                    when "0110100101000110" => rgb <= "010101";
                    when "0110100101000111" => rgb <= "010101";
                    when "0110100101001000" => rgb <= "010101";
                    when "0110100101001001" => rgb <= "010101";
                    when "0110100101001010" => rgb <= "010101";
                    when "0110100101001011" => rgb <= "010101";
                    when "0110100101001100" => rgb <= "010101";
                    when "0110100101001101" => rgb <= "010101";
                    when "0110100101001110" => rgb <= "010101";
                    when "0110100101010000" => rgb <= "101010";
                    when "0110100101010001" => rgb <= "101010";
                    when "0110100101010011" => rgb <= "010101";
                    when "0110100101010100" => rgb <= "010101";
                    when "0110100101010101" => rgb <= "101010";
                    when "0110100101011010" => rgb <= "101010";
                    when "0110100101011011" => rgb <= "101010";
                    when "0110100101011100" => rgb <= "010101";
                    when "0110100101011101" => rgb <= "010101";
                    when "0110100101011110" => rgb <= "010101";
                    when "0110100101011111" => rgb <= "010101";
                    when "0110100101100000" => rgb <= "010101";
                    when "0110100101100001" => rgb <= "010101";
                    when "0110100101100010" => rgb <= "010101";
                    when "0110100101100011" => rgb <= "010101";
                    when "0110100101100100" => rgb <= "010101";
                    when "0110100101100101" => rgb <= "010101";
                    when "0110100101100110" => rgb <= "010101";
                    when "0110100101100111" => rgb <= "010101";
                    when "0110100101101000" => rgb <= "010101";
                    when "0110100101101001" => rgb <= "010101";
                    when "0110100101101010" => rgb <= "010101";
                    when "0110100101101011" => rgb <= "010101";
                    when "0110100101101100" => rgb <= "010101";
                    when "0110100101101101" => rgb <= "010101";
                    when "0110100101101110" => rgb <= "010101";
                    when "0110100101101111" => rgb <= "010101";
                    when "0110100101110000" => rgb <= "101010";
                    when "0110100101110001" => rgb <= "101010";
                    when "0110100101110011" => rgb <= "010101";
                    when "0110100101110100" => rgb <= "010101";
                    when "0110100101110101" => rgb <= "010101";
                    when "0110100101110110" => rgb <= "010101";
                    when "0110100101110111" => rgb <= "010101";
                    when "0110100101111000" => rgb <= "010101";
                    when "0110100101111001" => rgb <= "010101";
                    when "0110100101111010" => rgb <= "010101";
                    when "0110100101111011" => rgb <= "010101";
                    when "0110100101111100" => rgb <= "010101";
                    when "0110100101111101" => rgb <= "010101";
                    when "0110100101111110" => rgb <= "010101";
                    when "0110100110000000" => rgb <= "101010";
                    when "0110100110000001" => rgb <= "101010";
                    when "0110100110000011" => rgb <= "010101";
                    when "0110100110000100" => rgb <= "010101";
                    when "0110100110000101" => rgb <= "010101";
                    when "0110100110000110" => rgb <= "010101";
                    when "0110100110010000" => rgb <= "101010";
                    when "0110100110010001" => rgb <= "101010";
                    when "0110100110010011" => rgb <= "010101";
                    when "0110100110010100" => rgb <= "010101";
                    when "0110100110010101" => rgb <= "010101";
                    when "0110100110010110" => rgb <= "010101";
                    when "0110100110010111" => rgb <= "010101";
                    when "0110100110011000" => rgb <= "010101";
                    when "0110100110011001" => rgb <= "010101";
                    when "0110100110011010" => rgb <= "010101";
                    when "0110100110011011" => rgb <= "010101";
                    when "0110100110011100" => rgb <= "010101";
                    when "0110100110011101" => rgb <= "010101";
                    when "0110100110011110" => rgb <= "010101";
                    when "0110101000000011" => rgb <= "010101";
                    when "0110101000000100" => rgb <= "010101";
                    when "0110101000000101" => rgb <= "010101";
                    when "0110101000000110" => rgb <= "010101";
                    when "0110101000000111" => rgb <= "010101";
                    when "0110101000001000" => rgb <= "010101";
                    when "0110101000001001" => rgb <= "010101";
                    when "0110101000001010" => rgb <= "010101";
                    when "0110101000001011" => rgb <= "010101";
                    when "0110101000001100" => rgb <= "010101";
                    when "0110101000001101" => rgb <= "010101";
                    when "0110101000001110" => rgb <= "010101";
                    when "0110101000010011" => rgb <= "010101";
                    when "0110101000010100" => rgb <= "010101";
                    when "0110101000101101" => rgb <= "010101";
                    when "0110101000101110" => rgb <= "010101";
                    when "0110101000110011" => rgb <= "010101";
                    when "0110101000110100" => rgb <= "010101";
                    when "0110101000110101" => rgb <= "010101";
                    when "0110101000110110" => rgb <= "010101";
                    when "0110101000110111" => rgb <= "010101";
                    when "0110101000111000" => rgb <= "010101";
                    when "0110101000111001" => rgb <= "010101";
                    when "0110101000111101" => rgb <= "010101";
                    when "0110101000111110" => rgb <= "010101";
                    when "0110101001000011" => rgb <= "010101";
                    when "0110101001001110" => rgb <= "010101";
                    when "0110101001010011" => rgb <= "010101";
                    when "0110101001010100" => rgb <= "010101";
                    when "0110101001010101" => rgb <= "101010";
                    when "0110101001011000" => rgb <= "101010";
                    when "0110101001011001" => rgb <= "101010";
                    when "0110101001011010" => rgb <= "010101";
                    when "0110101001011011" => rgb <= "010101";
                    when "0110101001011100" => rgb <= "010101";
                    when "0110101001011101" => rgb <= "010101";
                    when "0110101001011110" => rgb <= "010101";
                    when "0110101001011111" => rgb <= "010101";
                    when "0110101001100000" => rgb <= "010101";
                    when "0110101001100001" => rgb <= "010101";
                    when "0110101001100010" => rgb <= "010101";
                    when "0110101001100011" => rgb <= "010101";
                    when "0110101001100100" => rgb <= "010101";
                    when "0110101001100101" => rgb <= "010101";
                    when "0110101001100110" => rgb <= "010101";
                    when "0110101001100111" => rgb <= "010101";
                    when "0110101001101000" => rgb <= "010101";
                    when "0110101001101001" => rgb <= "010101";
                    when "0110101001101010" => rgb <= "010101";
                    when "0110101001101011" => rgb <= "010101";
                    when "0110101001101100" => rgb <= "010101";
                    when "0110101001101101" => rgb <= "010101";
                    when "0110101001101110" => rgb <= "010101";
                    when "0110101001101111" => rgb <= "010101";
                    when "0110101001110011" => rgb <= "010101";
                    when "0110101001110110" => rgb <= "010101";
                    when "0110101001110111" => rgb <= "010101";
                    when "0110101001111010" => rgb <= "010101";
                    when "0110101001111011" => rgb <= "010101";
                    when "0110101001111110" => rgb <= "010101";
                    when "0110101010000011" => rgb <= "010101";
                    when "0110101010000100" => rgb <= "010101";
                    when "0110101010000101" => rgb <= "010101";
                    when "0110101010000110" => rgb <= "010101";
                    when "0110101010000111" => rgb <= "010101";
                    when "0110101010001000" => rgb <= "010101";
                    when "0110101010001001" => rgb <= "010101";
                    when "0110101010001010" => rgb <= "010101";
                    when "0110101010001100" => rgb <= "010101";
                    when "0110101010001101" => rgb <= "010101";
                    when "0110101010001110" => rgb <= "010101";
                    when "0110101010010011" => rgb <= "010101";
                    when "0110101010010100" => rgb <= "010101";
                    when "0110101010010101" => rgb <= "010101";
                    when "0110101010010110" => rgb <= "010101";
                    when "0110101010010111" => rgb <= "010101";
                    when "0110101010011000" => rgb <= "010101";
                    when "0110101010011001" => rgb <= "010101";
                    when "0110101010011010" => rgb <= "010101";
                    when "0110101010011011" => rgb <= "010101";
                    when "0110101010011100" => rgb <= "010101";
                    when "0110101010011101" => rgb <= "010101";
                    when "0110101010011110" => rgb <= "010101";
                    when "0110101100000000" => rgb <= "101010";
                    when "0110101100000001" => rgb <= "101010";
                    when "0110101100000011" => rgb <= "010101";
                    when "0110101100000100" => rgb <= "010101";
                    when "0110101100001000" => rgb <= "010101";
                    when "0110101100001001" => rgb <= "010101";
                    when "0110101100001010" => rgb <= "010101";
                    when "0110101100001011" => rgb <= "010101";
                    when "0110101100001100" => rgb <= "010101";
                    when "0110101100001101" => rgb <= "010101";
                    when "0110101100001110" => rgb <= "010101";
                    when "0110101100010000" => rgb <= "101010";
                    when "0110101100010001" => rgb <= "101010";
                    when "0110101100010011" => rgb <= "010101";
                    when "0110101100010100" => rgb <= "010101";
                    when "0110101100010110" => rgb <= "010101";
                    when "0110101100010111" => rgb <= "010101";
                    when "0110101100011000" => rgb <= "010101";
                    when "0110101100011001" => rgb <= "010101";
                    when "0110101100011010" => rgb <= "010101";
                    when "0110101100011011" => rgb <= "010101";
                    when "0110101100011100" => rgb <= "010101";
                    when "0110101100011101" => rgb <= "010101";
                    when "0110101100011110" => rgb <= "010101";
                    when "0110101100100000" => rgb <= "101010";
                    when "0110101100100001" => rgb <= "101010";
                    when "0110101100100011" => rgb <= "010101";
                    when "0110101100100100" => rgb <= "010101";
                    when "0110101100100101" => rgb <= "010101";
                    when "0110101100100110" => rgb <= "010101";
                    when "0110101100100111" => rgb <= "010101";
                    when "0110101100101000" => rgb <= "010101";
                    when "0110101100101001" => rgb <= "010101";
                    when "0110101100101010" => rgb <= "010101";
                    when "0110101100101011" => rgb <= "010101";
                    when "0110101100101101" => rgb <= "010101";
                    when "0110101100101110" => rgb <= "010101";
                    when "0110101100110000" => rgb <= "101010";
                    when "0110101100110001" => rgb <= "101010";
                    when "0110101100110011" => rgb <= "010101";
                    when "0110101100110100" => rgb <= "010101";
                    when "0110101100110110" => rgb <= "010101";
                    when "0110101100111000" => rgb <= "010101";
                    when "0110101100111001" => rgb <= "010101";
                    when "0110101100111101" => rgb <= "010101";
                    when "0110101100111110" => rgb <= "010101";
                    when "0110101101000000" => rgb <= "101010";
                    when "0110101101000001" => rgb <= "101010";
                    when "0110101101000011" => rgb <= "010101";
                    when "0110101101001110" => rgb <= "010101";
                    when "0110101101010000" => rgb <= "101010";
                    when "0110101101010001" => rgb <= "101010";
                    when "0110101101010011" => rgb <= "010101";
                    when "0110101101010100" => rgb <= "010101";
                    when "0110101101010101" => rgb <= "101010";
                    when "0110101101011000" => rgb <= "010101";
                    when "0110101101011001" => rgb <= "010101";
                    when "0110101101011010" => rgb <= "010101";
                    when "0110101101011011" => rgb <= "010101";
                    when "0110101101011100" => rgb <= "010101";
                    when "0110101101011101" => rgb <= "010101";
                    when "0110101101100101" => rgb <= "010101";
                    when "0110101101100110" => rgb <= "010101";
                    when "0110101101100111" => rgb <= "010101";
                    when "0110101101101000" => rgb <= "010101";
                    when "0110101101101001" => rgb <= "010101";
                    when "0110101101101010" => rgb <= "010000";
                    when "0110101101101011" => rgb <= "010101";
                    when "0110101101101100" => rgb <= "010000";
                    when "0110101101101101" => rgb <= "010101";
                    when "0110101101101110" => rgb <= "010000";
                    when "0110101101101111" => rgb <= "010101";
                    when "0110101101110000" => rgb <= "101010";
                    when "0110101101110001" => rgb <= "101010";
                    when "0110101101110011" => rgb <= "010101";
                    when "0110101101110101" => rgb <= "010100";
                    when "0110101101110110" => rgb <= "010101";
                    when "0110101101110111" => rgb <= "010101";
                    when "0110101101111010" => rgb <= "010101";
                    when "0110101101111011" => rgb <= "010101";
                    when "0110101101111110" => rgb <= "010101";
                    when "0110101110000000" => rgb <= "101010";
                    when "0110101110000001" => rgb <= "101010";
                    when "0110101110000011" => rgb <= "010101";
                    when "0110101110000100" => rgb <= "010101";
                    when "0110101110001000" => rgb <= "010101";
                    when "0110101110001001" => rgb <= "010101";
                    when "0110101110001010" => rgb <= "010101";
                    when "0110101110001011" => rgb <= "010101";
                    when "0110101110001100" => rgb <= "010101";
                    when "0110101110001110" => rgb <= "010101";
                    when "0110101110010000" => rgb <= "101010";
                    when "0110101110010001" => rgb <= "101010";
                    when "0110101110010011" => rgb <= "010101";
                    when "0110101110010100" => rgb <= "010101";
                    when "0110101110010101" => rgb <= "010101";
                    when "0110101110010110" => rgb <= "010101";
                    when "0110101110010111" => rgb <= "010101";
                    when "0110101110011000" => rgb <= "010101";
                    when "0110101110011001" => rgb <= "010101";
                    when "0110101110011010" => rgb <= "010101";
                    when "0110101110011011" => rgb <= "010101";
                    when "0110101110011100" => rgb <= "010101";
                    when "0110101110011101" => rgb <= "010101";
                    when "0110101110011110" => rgb <= "010101";
                    when "0110110000000000" => rgb <= "101010";
                    when "0110110000000001" => rgb <= "101010";
                    when "0110110000000011" => rgb <= "010101";
                    when "0110110000000100" => rgb <= "010101";
                    when "0110110000001000" => rgb <= "010101";
                    when "0110110000001001" => rgb <= "010101";
                    when "0110110000001010" => rgb <= "010101";
                    when "0110110000001011" => rgb <= "010101";
                    when "0110110000001100" => rgb <= "010101";
                    when "0110110000001101" => rgb <= "010101";
                    when "0110110000001110" => rgb <= "010101";
                    when "0110110000010000" => rgb <= "101010";
                    when "0110110000010001" => rgb <= "101010";
                    when "0110110000010011" => rgb <= "010101";
                    when "0110110000010100" => rgb <= "010101";
                    when "0110110000010110" => rgb <= "010101";
                    when "0110110000010111" => rgb <= "010101";
                    when "0110110000011000" => rgb <= "101010";
                    when "0110110000011001" => rgb <= "010101";
                    when "0110110000011010" => rgb <= "101010";
                    when "0110110000011011" => rgb <= "101010";
                    when "0110110000011100" => rgb <= "010101";
                    when "0110110000011101" => rgb <= "101010";
                    when "0110110000011110" => rgb <= "101010";
                    when "0110110000100000" => rgb <= "101010";
                    when "0110110000100001" => rgb <= "101010";
                    when "0110110000100011" => rgb <= "101010";
                    when "0110110000100100" => rgb <= "101010";
                    when "0110110000100101" => rgb <= "010101";
                    when "0110110000100110" => rgb <= "101010";
                    when "0110110000100111" => rgb <= "101010";
                    when "0110110000101000" => rgb <= "010101";
                    when "0110110000101001" => rgb <= "101010";
                    when "0110110000101010" => rgb <= "010101";
                    when "0110110000101011" => rgb <= "010101";
                    when "0110110000101101" => rgb <= "010101";
                    when "0110110000101110" => rgb <= "010101";
                    when "0110110000110000" => rgb <= "101010";
                    when "0110110000110001" => rgb <= "101010";
                    when "0110110000110011" => rgb <= "010101";
                    when "0110110000110100" => rgb <= "010101";
                    when "0110110000110110" => rgb <= "010101";
                    when "0110110000111000" => rgb <= "010101";
                    when "0110110000111001" => rgb <= "010101";
                    when "0110110000111101" => rgb <= "010101";
                    when "0110110000111110" => rgb <= "010101";
                    when "0110110001000000" => rgb <= "101010";
                    when "0110110001000001" => rgb <= "101010";
                    when "0110110001000011" => rgb <= "010101";
                    when "0110110001001110" => rgb <= "010101";
                    when "0110110001010000" => rgb <= "101010";
                    when "0110110001010001" => rgb <= "101010";
                    when "0110110001010011" => rgb <= "010101";
                    when "0110110001010100" => rgb <= "010101";
                    when "0110110001010101" => rgb <= "101010";
                    when "0110110001011000" => rgb <= "010101";
                    when "0110110001011001" => rgb <= "010101";
                    when "0110110001011010" => rgb <= "010101";
                    when "0110110001011011" => rgb <= "010101";
                    when "0110110001100001" => rgb <= "010101";
                    when "0110110001100010" => rgb <= "010101";
                    when "0110110001100011" => rgb <= "010101";
                    when "0110110001100100" => rgb <= "010101";
                    when "0110110001100101" => rgb <= "010101";
                    when "0110110001100111" => rgb <= "010101";
                    when "0110110001101000" => rgb <= "010101";
                    when "0110110001101001" => rgb <= "010101";
                    when "0110110001101010" => rgb <= "010101";
                    when "0110110001101011" => rgb <= "010101";
                    when "0110110001101100" => rgb <= "010101";
                    when "0110110001101101" => rgb <= "010101";
                    when "0110110001101110" => rgb <= "010101";
                    when "0110110001101111" => rgb <= "010101";
                    when "0110110001110000" => rgb <= "101010";
                    when "0110110001110001" => rgb <= "101010";
                    when "0110110001110011" => rgb <= "010101";
                    when "0110110001110100" => rgb <= "010101";
                    when "0110110001110101" => rgb <= "010101";
                    when "0110110001110110" => rgb <= "010101";
                    when "0110110001110111" => rgb <= "010101";
                    when "0110110001111000" => rgb <= "010101";
                    when "0110110001111001" => rgb <= "010101";
                    when "0110110001111010" => rgb <= "010101";
                    when "0110110001111011" => rgb <= "010101";
                    when "0110110001111100" => rgb <= "010101";
                    when "0110110001111101" => rgb <= "010101";
                    when "0110110001111110" => rgb <= "010101";
                    when "0110110010000000" => rgb <= "101010";
                    when "0110110010000001" => rgb <= "101010";
                    when "0110110010000011" => rgb <= "010101";
                    when "0110110010000100" => rgb <= "010101";
                    when "0110110010001000" => rgb <= "010101";
                    when "0110110010001001" => rgb <= "010101";
                    when "0110110010001010" => rgb <= "010101";
                    when "0110110010001011" => rgb <= "010101";
                    when "0110110010001100" => rgb <= "010101";
                    when "0110110010001101" => rgb <= "010101";
                    when "0110110010001110" => rgb <= "010101";
                    when "0110110010010000" => rgb <= "101010";
                    when "0110110010010001" => rgb <= "101010";
                    when "0110110010010011" => rgb <= "010101";
                    when "0110110010010100" => rgb <= "010101";
                    when "0110110010011110" => rgb <= "010101";
                    when "0110110100000000" => rgb <= "101010";
                    when "0110110100000001" => rgb <= "101010";
                    when "0110110100000100" => rgb <= "010101";
                    when "0110110100001000" => rgb <= "010101";
                    when "0110110100001001" => rgb <= "010101";
                    when "0110110100001010" => rgb <= "010101";
                    when "0110110100001011" => rgb <= "010101";
                    when "0110110100001100" => rgb <= "010101";
                    when "0110110100001101" => rgb <= "010101";
                    when "0110110100001110" => rgb <= "010101";
                    when "0110110100010000" => rgb <= "101010";
                    when "0110110100010001" => rgb <= "101010";
                    when "0110110100010100" => rgb <= "010101";
                    when "0110110100010110" => rgb <= "010101";
                    when "0110110100010111" => rgb <= "101010";
                    when "0110110100011000" => rgb <= "000010";
                    when "0110110100011001" => rgb <= "010101";
                    when "0110110100011010" => rgb <= "100101";
                    when "0110110100011011" => rgb <= "000010";
                    when "0110110100011100" => rgb <= "010101";
                    when "0110110100011101" => rgb <= "000010";
                    when "0110110100011110" => rgb <= "000101";
                    when "0110110100100000" => rgb <= "101010";
                    when "0110110100100001" => rgb <= "101010";
                    when "0110110100100011" => rgb <= "000101";
                    when "0110110100100100" => rgb <= "000010";
                    when "0110110100100101" => rgb <= "010101";
                    when "0110110100100110" => rgb <= "000101";
                    when "0110110100100111" => rgb <= "000101";
                    when "0110110100101000" => rgb <= "010101";
                    when "0110110100101001" => rgb <= "100101";
                    when "0110110100101010" => rgb <= "101010";
                    when "0110110100101011" => rgb <= "010101";
                    when "0110110100101101" => rgb <= "010101";
                    when "0110110100101110" => rgb <= "010101";
                    when "0110110100110000" => rgb <= "101010";
                    when "0110110100110001" => rgb <= "101010";
                    when "0110110100110100" => rgb <= "010101";
                    when "0110110100110110" => rgb <= "010101";
                    when "0110110100111000" => rgb <= "010101";
                    when "0110110100111001" => rgb <= "010101";
                    when "0110110100111101" => rgb <= "010101";
                    when "0110110100111110" => rgb <= "010101";
                    when "0110110101000000" => rgb <= "101010";
                    when "0110110101000001" => rgb <= "101010";
                    when "0110110101000011" => rgb <= "010101";
                    when "0110110101001110" => rgb <= "010101";
                    when "0110110101010000" => rgb <= "101010";
                    when "0110110101010001" => rgb <= "101010";
                    when "0110110101010100" => rgb <= "010101";
                    when "0110110101010101" => rgb <= "101010";
                    when "0110110101010110" => rgb <= "101010";
                    when "0110110101010111" => rgb <= "010101";
                    when "0110110101011000" => rgb <= "010101";
                    when "0110110101011001" => rgb <= "010101";
                    when "0110110101011100" => rgb <= "010101";
                    when "0110110101011101" => rgb <= "010101";
                    when "0110110101011110" => rgb <= "101010";
                    when "0110110101011111" => rgb <= "101010";
                    when "0110110101100000" => rgb <= "101010";
                    when "0110110101100001" => rgb <= "101010";
                    when "0110110101100010" => rgb <= "010101";
                    when "0110110101100011" => rgb <= "010101";
                    when "0110110101100100" => rgb <= "010101";
                    when "0110110101100101" => rgb <= "010101";
                    when "0110110101100110" => rgb <= "010101";
                    when "0110110101100111" => rgb <= "010101";
                    when "0110110101101001" => rgb <= "010101";
                    when "0110110101101010" => rgb <= "010101";
                    when "0110110101101011" => rgb <= "010101";
                    when "0110110101101100" => rgb <= "010101";
                    when "0110110101101101" => rgb <= "010101";
                    when "0110110101101110" => rgb <= "010000";
                    when "0110110101101111" => rgb <= "010101";
                    when "0110110101110000" => rgb <= "101010";
                    when "0110110101110001" => rgb <= "101010";
                    when "0110110101110011" => rgb <= "010101";
                    when "0110110101110100" => rgb <= "010101";
                    when "0110110101110101" => rgb <= "010101";
                    when "0110110101110110" => rgb <= "010101";
                    when "0110110101110111" => rgb <= "010101";
                    when "0110110101111000" => rgb <= "010101";
                    when "0110110101111001" => rgb <= "010101";
                    when "0110110101111010" => rgb <= "010101";
                    when "0110110101111011" => rgb <= "010101";
                    when "0110110101111100" => rgb <= "010101";
                    when "0110110101111101" => rgb <= "010101";
                    when "0110110101111110" => rgb <= "010101";
                    when "0110110110000000" => rgb <= "101010";
                    when "0110110110000001" => rgb <= "101010";
                    when "0110110110000100" => rgb <= "010101";
                    when "0110110110001000" => rgb <= "010101";
                    when "0110110110001001" => rgb <= "010101";
                    when "0110110110001010" => rgb <= "010101";
                    when "0110110110001011" => rgb <= "010101";
                    when "0110110110001100" => rgb <= "010101";
                    when "0110110110001101" => rgb <= "010101";
                    when "0110110110001110" => rgb <= "010101";
                    when "0110110110010000" => rgb <= "101010";
                    when "0110110110010001" => rgb <= "101010";
                    when "0110110110010100" => rgb <= "010101";
                    when "0110110110011110" => rgb <= "010101";
                    when "0110111000000100" => rgb <= "010101";
                    when "0110111000001000" => rgb <= "010101";
                    when "0110111000001001" => rgb <= "010101";
                    when "0110111000001010" => rgb <= "010101";
                    when "0110111000001011" => rgb <= "010101";
                    when "0110111000001100" => rgb <= "010101";
                    when "0110111000001101" => rgb <= "010101";
                    when "0110111000001110" => rgb <= "010101";
                    when "0110111000010100" => rgb <= "010101";
                    when "0110111000010110" => rgb <= "010101";
                    when "0110111000010111" => rgb <= "000010";
                    when "0110111000011000" => rgb <= "000010";
                    when "0110111000011001" => rgb <= "010101";
                    when "0110111000011010" => rgb <= "000010";
                    when "0110111000011011" => rgb <= "000010";
                    when "0110111000011100" => rgb <= "010101";
                    when "0110111000011101" => rgb <= "000101";
                    when "0110111000011110" => rgb <= "000010";
                    when "0110111000100011" => rgb <= "100101";
                    when "0110111000100100" => rgb <= "000010";
                    when "0110111000100101" => rgb <= "010101";
                    when "0110111000100110" => rgb <= "100101";
                    when "0110111000100111" => rgb <= "000101";
                    when "0110111000101000" => rgb <= "010101";
                    when "0110111000101001" => rgb <= "000101";
                    when "0110111000101010" => rgb <= "100101";
                    when "0110111000101011" => rgb <= "010101";
                    when "0110111000101101" => rgb <= "010101";
                    when "0110111000101110" => rgb <= "010101";
                    when "0110111000110100" => rgb <= "010101";
                    when "0110111000110110" => rgb <= "010101";
                    when "0110111000111000" => rgb <= "010101";
                    when "0110111000111001" => rgb <= "010101";
                    when "0110111000111101" => rgb <= "010101";
                    when "0110111000111110" => rgb <= "010101";
                    when "0110111001000011" => rgb <= "010101";
                    when "0110111001001110" => rgb <= "010101";
                    when "0110111001010100" => rgb <= "010101";
                    when "0110111001010101" => rgb <= "101010";
                    when "0110111001010110" => rgb <= "010101";
                    when "0110111001010111" => rgb <= "010101";
                    when "0110111001011000" => rgb <= "010101";
                    when "0110111001011010" => rgb <= "010101";
                    when "0110111001011011" => rgb <= "010101";
                    when "0110111001011100" => rgb <= "101010";
                    when "0110111001011101" => rgb <= "010101";
                    when "0110111001011110" => rgb <= "010101";
                    when "0110111001011111" => rgb <= "010101";
                    when "0110111001100000" => rgb <= "010101";
                    when "0110111001100001" => rgb <= "010101";
                    when "0110111001100010" => rgb <= "010101";
                    when "0110111001100011" => rgb <= "010101";
                    when "0110111001100100" => rgb <= "010101";
                    when "0110111001100101" => rgb <= "010101";
                    when "0110111001100110" => rgb <= "010101";
                    when "0110111001100111" => rgb <= "010101";
                    when "0110111001101000" => rgb <= "010101";
                    when "0110111001101010" => rgb <= "010101";
                    when "0110111001101011" => rgb <= "010101";
                    when "0110111001101100" => rgb <= "010101";
                    when "0110111001101101" => rgb <= "010101";
                    when "0110111001101110" => rgb <= "010101";
                    when "0110111001101111" => rgb <= "010101";
                    when "0110111001110011" => rgb <= "010101";
                    when "0110111001110110" => rgb <= "010101";
                    when "0110111001110111" => rgb <= "010101";
                    when "0110111001111010" => rgb <= "010101";
                    when "0110111001111011" => rgb <= "010101";
                    when "0110111001111101" => rgb <= "100000";
                    when "0110111001111110" => rgb <= "010101";
                    when "0110111010000100" => rgb <= "010101";
                    when "0110111010001000" => rgb <= "010101";
                    when "0110111010001001" => rgb <= "010101";
                    when "0110111010001100" => rgb <= "010101";
                    when "0110111010001101" => rgb <= "010101";
                    when "0110111010001110" => rgb <= "010101";
                    when "0110111010010100" => rgb <= "010101";
                    when "0110111010010110" => rgb <= "100000";
                    when "0110111010010111" => rgb <= "000010";
                    when "0110111010011000" => rgb <= "100101";
                    when "0110111010011001" => rgb <= "010100";
                    when "0110111010011010" => rgb <= "000010";
                    when "0110111010011011" => rgb <= "010100";
                    when "0110111010011100" => rgb <= "100000";
                    when "0110111010011110" => rgb <= "010101";
                    when "0110111100000100" => rgb <= "010101";
                    when "0110111100001000" => rgb <= "010101";
                    when "0110111100001001" => rgb <= "010101";
                    when "0110111100001010" => rgb <= "010101";
                    when "0110111100001011" => rgb <= "010101";
                    when "0110111100001100" => rgb <= "010101";
                    when "0110111100001101" => rgb <= "010101";
                    when "0110111100001110" => rgb <= "010101";
                    when "0110111100010100" => rgb <= "010101";
                    when "0110111100010110" => rgb <= "010101";
                    when "0110111100010111" => rgb <= "100101";
                    when "0110111100011000" => rgb <= "000101";
                    when "0110111100011001" => rgb <= "010101";
                    when "0110111100011010" => rgb <= "000010";
                    when "0110111100011011" => rgb <= "000101";
                    when "0110111100011100" => rgb <= "010101";
                    when "0110111100011101" => rgb <= "000010";
                    when "0110111100011110" => rgb <= "100101";
                    when "0110111100100011" => rgb <= "100101";
                    when "0110111100100100" => rgb <= "000101";
                    when "0110111100100101" => rgb <= "010101";
                    when "0110111100100110" => rgb <= "000010";
                    when "0110111100100111" => rgb <= "100101";
                    when "0110111100101000" => rgb <= "010101";
                    when "0110111100101001" => rgb <= "000101";
                    when "0110111100101010" => rgb <= "000010";
                    when "0110111100101011" => rgb <= "010101";
                    when "0110111100101101" => rgb <= "010101";
                    when "0110111100101110" => rgb <= "010101";
                    when "0110111100110100" => rgb <= "010101";
                    when "0110111100110110" => rgb <= "010101";
                    when "0110111100111000" => rgb <= "010101";
                    when "0110111100111001" => rgb <= "010101";
                    when "0110111100111010" => rgb <= "010101";
                    when "0110111100111011" => rgb <= "010101";
                    when "0110111100111100" => rgb <= "010101";
                    when "0110111100111101" => rgb <= "010101";
                    when "0110111100111110" => rgb <= "010101";
                    when "0110111101000011" => rgb <= "010101";
                    when "0110111101000100" => rgb <= "010101";
                    when "0110111101000101" => rgb <= "010101";
                    when "0110111101000110" => rgb <= "010101";
                    when "0110111101000111" => rgb <= "010101";
                    when "0110111101001000" => rgb <= "010101";
                    when "0110111101001001" => rgb <= "010101";
                    when "0110111101001010" => rgb <= "010101";
                    when "0110111101001011" => rgb <= "010101";
                    when "0110111101001100" => rgb <= "010101";
                    when "0110111101001101" => rgb <= "010101";
                    when "0110111101001110" => rgb <= "010101";
                    when "0110111101010100" => rgb <= "010101";
                    when "0110111101010101" => rgb <= "101010";
                    when "0110111101010110" => rgb <= "010101";
                    when "0110111101010111" => rgb <= "010101";
                    when "0110111101011010" => rgb <= "010101";
                    when "0110111101011011" => rgb <= "010101";
                    when "0110111101011100" => rgb <= "010101";
                    when "0110111101011101" => rgb <= "010101";
                    when "0110111101011110" => rgb <= "010101";
                    when "0110111101011111" => rgb <= "010101";
                    when "0110111101100000" => rgb <= "010101";
                    when "0110111101100001" => rgb <= "010101";
                    when "0110111101100010" => rgb <= "010101";
                    when "0110111101100011" => rgb <= "010101";
                    when "0110111101100100" => rgb <= "010101";
                    when "0110111101100101" => rgb <= "010101";
                    when "0110111101100110" => rgb <= "010101";
                    when "0110111101100111" => rgb <= "010101";
                    when "0110111101101000" => rgb <= "010101";
                    when "0110111101101001" => rgb <= "010101";
                    when "0110111101101011" => rgb <= "010101";
                    when "0110111101101100" => rgb <= "010101";
                    when "0110111101101101" => rgb <= "010101";
                    when "0110111101101110" => rgb <= "010000";
                    when "0110111101101111" => rgb <= "010101";
                    when "0110111101110011" => rgb <= "010101";
                    when "0110111101110100" => rgb <= "100000";
                    when "0110111101110110" => rgb <= "010101";
                    when "0110111101110111" => rgb <= "010101";
                    when "0110111101111010" => rgb <= "010101";
                    when "0110111101111011" => rgb <= "010101";
                    when "0110111101111110" => rgb <= "010101";
                    when "0110111110000100" => rgb <= "010101";
                    when "0110111110001000" => rgb <= "010101";
                    when "0110111110001001" => rgb <= "010101";
                    when "0110111110001100" => rgb <= "010101";
                    when "0110111110001101" => rgb <= "010101";
                    when "0110111110001110" => rgb <= "010101";
                    when "0110111110010100" => rgb <= "010101";
                    when "0110111110010110" => rgb <= "000010";
                    when "0110111110010111" => rgb <= "100000";
                    when "0110111110011000" => rgb <= "000010";
                    when "0110111110011001" => rgb <= "100000";
                    when "0110111110011010" => rgb <= "010100";
                    when "0110111110011011" => rgb <= "000010";
                    when "0110111110011100" => rgb <= "000010";
                    when "0110111110011110" => rgb <= "010101";
                    when "0111000000000000" => rgb <= "101010";
                    when "0111000000000001" => rgb <= "101010";
                    when "0111000000000100" => rgb <= "010101";
                    when "0111000000000101" => rgb <= "010101";
                    when "0111000000000110" => rgb <= "010101";
                    when "0111000000000111" => rgb <= "010101";
                    when "0111000000001000" => rgb <= "010101";
                    when "0111000000001001" => rgb <= "010101";
                    when "0111000000001101" => rgb <= "010101";
                    when "0111000000001110" => rgb <= "010101";
                    when "0111000000010000" => rgb <= "101010";
                    when "0111000000010001" => rgb <= "101010";
                    when "0111000000010100" => rgb <= "010101";
                    when "0111000000010110" => rgb <= "010101";
                    when "0111000000010111" => rgb <= "101010";
                    when "0111000000011000" => rgb <= "101010";
                    when "0111000000011001" => rgb <= "010101";
                    when "0111000000011010" => rgb <= "101010";
                    when "0111000000011011" => rgb <= "101010";
                    when "0111000000011100" => rgb <= "010101";
                    when "0111000000011101" => rgb <= "101010";
                    when "0111000000011110" => rgb <= "101010";
                    when "0111000000100000" => rgb <= "101010";
                    when "0111000000100001" => rgb <= "101010";
                    when "0111000000100011" => rgb <= "101010";
                    when "0111000000100100" => rgb <= "101010";
                    when "0111000000100101" => rgb <= "010101";
                    when "0111000000100110" => rgb <= "101010";
                    when "0111000000100111" => rgb <= "101010";
                    when "0111000000101000" => rgb <= "010101";
                    when "0111000000101001" => rgb <= "101010";
                    when "0111000000101010" => rgb <= "101010";
                    when "0111000000101011" => rgb <= "010101";
                    when "0111000000101101" => rgb <= "010101";
                    when "0111000000101110" => rgb <= "010101";
                    when "0111000000110000" => rgb <= "101010";
                    when "0111000000110001" => rgb <= "101010";
                    when "0111000000110100" => rgb <= "010101";
                    when "0111000000110101" => rgb <= "010101";
                    when "0111000000110110" => rgb <= "010101";
                    when "0111000000110111" => rgb <= "010101";
                    when "0111000000111000" => rgb <= "010101";
                    when "0111000000111001" => rgb <= "010101";
                    when "0111000000111010" => rgb <= "010101";
                    when "0111000000111011" => rgb <= "010101";
                    when "0111000000111100" => rgb <= "010101";
                    when "0111000000111101" => rgb <= "010101";
                    when "0111000000111110" => rgb <= "010101";
                    when "0111000001000000" => rgb <= "101010";
                    when "0111000001000001" => rgb <= "101010";
                    when "0111000001000100" => rgb <= "010101";
                    when "0111000001001110" => rgb <= "010101";
                    when "0111000001010000" => rgb <= "101010";
                    when "0111000001010001" => rgb <= "101010";
                    when "0111000001010100" => rgb <= "010101";
                    when "0111000001010101" => rgb <= "010101";
                    when "0111000001010110" => rgb <= "010101";
                    when "0111000001010111" => rgb <= "010101";
                    when "0111000001011001" => rgb <= "010101";
                    when "0111000001011010" => rgb <= "101010";
                    when "0111000001011011" => rgb <= "010101";
                    when "0111000001011100" => rgb <= "010101";
                    when "0111000001011101" => rgb <= "010101";
                    when "0111000001011110" => rgb <= "010101";
                    when "0111000001011111" => rgb <= "010101";
                    when "0111000001100000" => rgb <= "010101";
                    when "0111000001100001" => rgb <= "010101";
                    when "0111000001100010" => rgb <= "010101";
                    when "0111000001100011" => rgb <= "010101";
                    when "0111000001100100" => rgb <= "010101";
                    when "0111000001100101" => rgb <= "010101";
                    when "0111000001100110" => rgb <= "010101";
                    when "0111000001100111" => rgb <= "010101";
                    when "0111000001101000" => rgb <= "010101";
                    when "0111000001101001" => rgb <= "010101";
                    when "0111000001101011" => rgb <= "010101";
                    when "0111000001101100" => rgb <= "010101";
                    when "0111000001101101" => rgb <= "010101";
                    when "0111000001101110" => rgb <= "010101";
                    when "0111000001101111" => rgb <= "010101";
                    when "0111000001110000" => rgb <= "101010";
                    when "0111000001110001" => rgb <= "101010";
                    when "0111000001110011" => rgb <= "010101";
                    when "0111000001110100" => rgb <= "010101";
                    when "0111000001110101" => rgb <= "010101";
                    when "0111000001110110" => rgb <= "010101";
                    when "0111000001110111" => rgb <= "010101";
                    when "0111000001111000" => rgb <= "010101";
                    when "0111000001111001" => rgb <= "010101";
                    when "0111000001111010" => rgb <= "010101";
                    when "0111000001111011" => rgb <= "010101";
                    when "0111000001111100" => rgb <= "010101";
                    when "0111000001111101" => rgb <= "010101";
                    when "0111000001111110" => rgb <= "010101";
                    when "0111000010000000" => rgb <= "101010";
                    when "0111000010000001" => rgb <= "101010";
                    when "0111000010000100" => rgb <= "010101";
                    when "0111000010000101" => rgb <= "010101";
                    when "0111000010000110" => rgb <= "010101";
                    when "0111000010000111" => rgb <= "010101";
                    when "0111000010001000" => rgb <= "010101";
                    when "0111000010001001" => rgb <= "010101";
                    when "0111000010001100" => rgb <= "010101";
                    when "0111000010001101" => rgb <= "010101";
                    when "0111000010001110" => rgb <= "010101";
                    when "0111000010010000" => rgb <= "101010";
                    when "0111000010010001" => rgb <= "101010";
                    when "0111000010010100" => rgb <= "010101";
                    when "0111000010011110" => rgb <= "010101";
                    when "0111000100000000" => rgb <= "101010";
                    when "0111000100000001" => rgb <= "101010";
                    when "0111000100000100" => rgb <= "010101";
                    when "0111000100000101" => rgb <= "010101";
                    when "0111000100000110" => rgb <= "010101";
                    when "0111000100000111" => rgb <= "010101";
                    when "0111000100001000" => rgb <= "010101";
                    when "0111000100001001" => rgb <= "010101";
                    when "0111000100001101" => rgb <= "010101";
                    when "0111000100010000" => rgb <= "101010";
                    when "0111000100010001" => rgb <= "101010";
                    when "0111000100010100" => rgb <= "010101";
                    when "0111000100010110" => rgb <= "010101";
                    when "0111000100010111" => rgb <= "010101";
                    when "0111000100011000" => rgb <= "010101";
                    when "0111000100011001" => rgb <= "010101";
                    when "0111000100011010" => rgb <= "010101";
                    when "0111000100011011" => rgb <= "010101";
                    when "0111000100011100" => rgb <= "010101";
                    when "0111000100011101" => rgb <= "010101";
                    when "0111000100100000" => rgb <= "101010";
                    when "0111000100100001" => rgb <= "101010";
                    when "0111000100100100" => rgb <= "010101";
                    when "0111000100100101" => rgb <= "010101";
                    when "0111000100100110" => rgb <= "010101";
                    when "0111000100100111" => rgb <= "010101";
                    when "0111000100101000" => rgb <= "010101";
                    when "0111000100101001" => rgb <= "010101";
                    when "0111000100101010" => rgb <= "010101";
                    when "0111000100101011" => rgb <= "010101";
                    when "0111000100101101" => rgb <= "010101";
                    when "0111000100110000" => rgb <= "101010";
                    when "0111000100110001" => rgb <= "101010";
                    when "0111000100110100" => rgb <= "010101";
                    when "0111000100110111" => rgb <= "010101";
                    when "0111000100111000" => rgb <= "010101";
                    when "0111000100111100" => rgb <= "010101";
                    when "0111000100111101" => rgb <= "010101";
                    when "0111000101000000" => rgb <= "101010";
                    when "0111000101000001" => rgb <= "101010";
                    when "0111000101000100" => rgb <= "010101";
                    when "0111000101000111" => rgb <= "101010";
                    when "0111000101001001" => rgb <= "101010";
                    when "0111000101001011" => rgb <= "101010";
                    when "0111000101001110" => rgb <= "010101";
                    when "0111000101010000" => rgb <= "101010";
                    when "0111000101010001" => rgb <= "101010";
                    when "0111000101010100" => rgb <= "010101";
                    when "0111000101010101" => rgb <= "010101";
                    when "0111000101010110" => rgb <= "010101";
                    when "0111000101011000" => rgb <= "010101";
                    when "0111000101011001" => rgb <= "101010";
                    when "0111000101011010" => rgb <= "010101";
                    when "0111000101011011" => rgb <= "010101";
                    when "0111000101011100" => rgb <= "010101";
                    when "0111000101011101" => rgb <= "010101";
                    when "0111000101011110" => rgb <= "010101";
                    when "0111000101011111" => rgb <= "010101";
                    when "0111000101100000" => rgb <= "010101";
                    when "0111000101100001" => rgb <= "010101";
                    when "0111000101100010" => rgb <= "010101";
                    when "0111000101100011" => rgb <= "010101";
                    when "0111000101100100" => rgb <= "010101";
                    when "0111000101100101" => rgb <= "010101";
                    when "0111000101100110" => rgb <= "010101";
                    when "0111000101100111" => rgb <= "010101";
                    when "0111000101101000" => rgb <= "010101";
                    when "0111000101101001" => rgb <= "101010";
                    when "0111000101101010" => rgb <= "010101";
                    when "0111000101101100" => rgb <= "010101";
                    when "0111000101101101" => rgb <= "010101";
                    when "0111000101101110" => rgb <= "010101";
                    when "0111000101101111" => rgb <= "010101";
                    when "0111000101110000" => rgb <= "101010";
                    when "0111000101110001" => rgb <= "101010";
                    when "0111000101110011" => rgb <= "010101";
                    when "0111000101110100" => rgb <= "010101";
                    when "0111000101110101" => rgb <= "010101";
                    when "0111000101110110" => rgb <= "010101";
                    when "0111000101110111" => rgb <= "010101";
                    when "0111000101111000" => rgb <= "010101";
                    when "0111000101111001" => rgb <= "010101";
                    when "0111000101111010" => rgb <= "010101";
                    when "0111000101111011" => rgb <= "010101";
                    when "0111000101111100" => rgb <= "010101";
                    when "0111000101111101" => rgb <= "010101";
                    when "0111000101111110" => rgb <= "010101";
                    when "0111000110000000" => rgb <= "101010";
                    when "0111000110000001" => rgb <= "101010";
                    when "0111000110000100" => rgb <= "010101";
                    when "0111000110000111" => rgb <= "010101";
                    when "0111000110001000" => rgb <= "010101";
                    when "0111000110001001" => rgb <= "010101";
                    when "0111000110001010" => rgb <= "010101";
                    when "0111000110001011" => rgb <= "010101";
                    when "0111000110001100" => rgb <= "010101";
                    when "0111000110001101" => rgb <= "010101";
                    when "0111000110010000" => rgb <= "101010";
                    when "0111000110010001" => rgb <= "101010";
                    when "0111000110010100" => rgb <= "010101";
                    when "0111000110011110" => rgb <= "010101";
                    when "0111001000000100" => rgb <= "010101";
                    when "0111001000000101" => rgb <= "010101";
                    when "0111001000000110" => rgb <= "010101";
                    when "0111001000000111" => rgb <= "010101";
                    when "0111001000001000" => rgb <= "010101";
                    when "0111001000001001" => rgb <= "010101";
                    when "0111001000001101" => rgb <= "010101";
                    when "0111001000010100" => rgb <= "010101";
                    when "0111001000101101" => rgb <= "010101";
                    when "0111001000110100" => rgb <= "010101";
                    when "0111001000110101" => rgb <= "010101";
                    when "0111001000110111" => rgb <= "010101";
                    when "0111001000111000" => rgb <= "010101";
                    when "0111001000111100" => rgb <= "010101";
                    when "0111001000111101" => rgb <= "010101";
                    when "0111001001000011" => rgb <= "010101";
                    when "0111001001000100" => rgb <= "010101";
                    when "0111001001000101" => rgb <= "101010";
                    when "0111001001000110" => rgb <= "010101";
                    when "0111001001000111" => rgb <= "010101";
                    when "0111001001001000" => rgb <= "010101";
                    when "0111001001001001" => rgb <= "010101";
                    when "0111001001001010" => rgb <= "010101";
                    when "0111001001001011" => rgb <= "010101";
                    when "0111001001001100" => rgb <= "010101";
                    when "0111001001001101" => rgb <= "101010";
                    when "0111001001010100" => rgb <= "010101";
                    when "0111001001010101" => rgb <= "010101";
                    when "0111001001010110" => rgb <= "010101";
                    when "0111001001010111" => rgb <= "010101";
                    when "0111001001011000" => rgb <= "010101";
                    when "0111001001011001" => rgb <= "010101";
                    when "0111001001011010" => rgb <= "010101";
                    when "0111001001011011" => rgb <= "010101";
                    when "0111001001011100" => rgb <= "010101";
                    when "0111001001011101" => rgb <= "010101";
                    when "0111001001011110" => rgb <= "010101";
                    when "0111001001011111" => rgb <= "010101";
                    when "0111001001100000" => rgb <= "010101";
                    when "0111001001100001" => rgb <= "010101";
                    when "0111001001100010" => rgb <= "010101";
                    when "0111001001100011" => rgb <= "010101";
                    when "0111001001100100" => rgb <= "010101";
                    when "0111001001100101" => rgb <= "010101";
                    when "0111001001100110" => rgb <= "010101";
                    when "0111001001100111" => rgb <= "010101";
                    when "0111001001101000" => rgb <= "010101";
                    when "0111001001101001" => rgb <= "010101";
                    when "0111001001101010" => rgb <= "010101";
                    when "0111001001101011" => rgb <= "010101";
                    when "0111001001101100" => rgb <= "010101";
                    when "0111001001101101" => rgb <= "010101";
                    when "0111001001101111" => rgb <= "010101";
                    when "0111001001110011" => rgb <= "010101";
                    when "0111001001110110" => rgb <= "010101";
                    when "0111001001110111" => rgb <= "010101";
                    when "0111001001111010" => rgb <= "010101";
                    when "0111001001111011" => rgb <= "010101";
                    when "0111001001111100" => rgb <= "100000";
                    when "0111001001111110" => rgb <= "010101";
                    when "0111001010000100" => rgb <= "010101";
                    when "0111001010001000" => rgb <= "010101";
                    when "0111001010001001" => rgb <= "010101";
                    when "0111001010001100" => rgb <= "010101";
                    when "0111001010001101" => rgb <= "010101";
                    when "0111001010010100" => rgb <= "010101";
                    when "0111001010010101" => rgb <= "010101";
                    when "0111001010010111" => rgb <= "010101";
                    when "0111001010011000" => rgb <= "010101";
                    when "0111001010011001" => rgb <= "010101";
                    when "0111001010011110" => rgb <= "010101";
                    when "0111001100000100" => rgb <= "010101";
                    when "0111001100000101" => rgb <= "010101";
                    when "0111001100000110" => rgb <= "010101";
                    when "0111001100000111" => rgb <= "010101";
                    when "0111001100001000" => rgb <= "010101";
                    when "0111001100001001" => rgb <= "010101";
                    when "0111001100001100" => rgb <= "010101";
                    when "0111001100001101" => rgb <= "010101";
                    when "0111001100010100" => rgb <= "010101";
                    when "0111001100010101" => rgb <= "010101";
                    when "0111001100010110" => rgb <= "010101";
                    when "0111001100010111" => rgb <= "010101";
                    when "0111001100011000" => rgb <= "010101";
                    when "0111001100011001" => rgb <= "010101";
                    when "0111001100011010" => rgb <= "010101";
                    when "0111001100011011" => rgb <= "010101";
                    when "0111001100011100" => rgb <= "010101";
                    when "0111001100011101" => rgb <= "010101";
                    when "0111001100100100" => rgb <= "010101";
                    when "0111001100100101" => rgb <= "010101";
                    when "0111001100100110" => rgb <= "010101";
                    when "0111001100100111" => rgb <= "010101";
                    when "0111001100101000" => rgb <= "010101";
                    when "0111001100101001" => rgb <= "010101";
                    when "0111001100101010" => rgb <= "010101";
                    when "0111001100101011" => rgb <= "010101";
                    when "0111001100101100" => rgb <= "010101";
                    when "0111001100101101" => rgb <= "010101";
                    when "0111001100110100" => rgb <= "010101";
                    when "0111001100110101" => rgb <= "010101";
                    when "0111001100110110" => rgb <= "010101";
                    when "0111001100110111" => rgb <= "010101";
                    when "0111001100111000" => rgb <= "010101";
                    when "0111001100111001" => rgb <= "010101";
                    when "0111001100111100" => rgb <= "010101";
                    when "0111001100111101" => rgb <= "010101";
                    when "0111001101000100" => rgb <= "010101";
                    when "0111001101000101" => rgb <= "010101";
                    when "0111001101000111" => rgb <= "010101";
                    when "0111001101001000" => rgb <= "010101";
                    when "0111001101001001" => rgb <= "010101";
                    when "0111001101001011" => rgb <= "010101";
                    when "0111001101001100" => rgb <= "010101";
                    when "0111001101001101" => rgb <= "010101";
                    when "0111001101010100" => rgb <= "010101";
                    when "0111001101010101" => rgb <= "010101";
                    when "0111001101010111" => rgb <= "010101";
                    when "0111001101011000" => rgb <= "010101";
                    when "0111001101011001" => rgb <= "010101";
                    when "0111001101011010" => rgb <= "010101";
                    when "0111001101011011" => rgb <= "010101";
                    when "0111001101011100" => rgb <= "010101";
                    when "0111001101011101" => rgb <= "010101";
                    when "0111001101011110" => rgb <= "010101";
                    when "0111001101011111" => rgb <= "010101";
                    when "0111001101100000" => rgb <= "010101";
                    when "0111001101100001" => rgb <= "010101";
                    when "0111001101100010" => rgb <= "010101";
                    when "0111001101100011" => rgb <= "010101";
                    when "0111001101100100" => rgb <= "010101";
                    when "0111001101100101" => rgb <= "010101";
                    when "0111001101100110" => rgb <= "010101";
                    when "0111001101100111" => rgb <= "010101";
                    when "0111001101101000" => rgb <= "010101";
                    when "0111001101101001" => rgb <= "010101";
                    when "0111001101101010" => rgb <= "010101";
                    when "0111001101101011" => rgb <= "010101";
                    when "0111001101101101" => rgb <= "010101";
                    when "0111001101101111" => rgb <= "010101";
                    when "0111001101110011" => rgb <= "010101";
                    when "0111001101110110" => rgb <= "010101";
                    when "0111001101110111" => rgb <= "010101";
                    when "0111001101111000" => rgb <= "010100";
                    when "0111001101111010" => rgb <= "010101";
                    when "0111001101111011" => rgb <= "010101";
                    when "0111001101111101" => rgb <= "010100";
                    when "0111001101111110" => rgb <= "010101";
                    when "0111001110000100" => rgb <= "010101";
                    when "0111001110000101" => rgb <= "010101";
                    when "0111001110000110" => rgb <= "010101";
                    when "0111001110000111" => rgb <= "010101";
                    when "0111001110001000" => rgb <= "010101";
                    when "0111001110001001" => rgb <= "010101";
                    when "0111001110001100" => rgb <= "010101";
                    when "0111001110001101" => rgb <= "010101";
                    when "0111001110001110" => rgb <= "010101";
                    when "0111001110010100" => rgb <= "010101";
                    when "0111001110010101" => rgb <= "010101";
                    when "0111001110010110" => rgb <= "010101";
                    when "0111001110010111" => rgb <= "010101";
                    when "0111001110011000" => rgb <= "010101";
                    when "0111001110011001" => rgb <= "010101";
                    when "0111001110011010" => rgb <= "010101";
                    when "0111001110011011" => rgb <= "010101";
                    when "0111001110011100" => rgb <= "010101";
                    when "0111001110011101" => rgb <= "010101";
                    when "0111001110011110" => rgb <= "010101";
                    when "0111010000000100" => rgb <= "010101";
                    when "0111010000000101" => rgb <= "010101";
                    when "0111010000000110" => rgb <= "010101";
                    when "0111010000000111" => rgb <= "010101";
                    when "0111010000001001" => rgb <= "010101";
                    when "0111010000001100" => rgb <= "010101";
                    when "0111010000010100" => rgb <= "010101";
                    when "0111010000010111" => rgb <= "010101";
                    when "0111010000011001" => rgb <= "010101";
                    when "0111010000011010" => rgb <= "010101";
                    when "0111010000011100" => rgb <= "010101";
                    when "0111010000100100" => rgb <= "010101";
                    when "0111010000100101" => rgb <= "010101";
                    when "0111010000100110" => rgb <= "010101";
                    when "0111010000100111" => rgb <= "010101";
                    when "0111010000101001" => rgb <= "010101";
                    when "0111010000101010" => rgb <= "010101";
                    when "0111010000101011" => rgb <= "010101";
                    when "0111010000101100" => rgb <= "010101";
                    when "0111010000110100" => rgb <= "010101";
                    when "0111010000110101" => rgb <= "010101";
                    when "0111010000110110" => rgb <= "010101";
                    when "0111010000110111" => rgb <= "010101";
                    when "0111010000111001" => rgb <= "010101";
                    when "0111010000111100" => rgb <= "010101";
                    when "0111010001000100" => rgb <= "010101";
                    when "0111010001000101" => rgb <= "010101";
                    when "0111010001000110" => rgb <= "010101";
                    when "0111010001000111" => rgb <= "010101";
                    when "0111010001001000" => rgb <= "010101";
                    when "0111010001001001" => rgb <= "010101";
                    when "0111010001001010" => rgb <= "010101";
                    when "0111010001001011" => rgb <= "010101";
                    when "0111010001001100" => rgb <= "010101";
                    when "0111010001001101" => rgb <= "010101";
                    when "0111010001010100" => rgb <= "010101";
                    when "0111010001010101" => rgb <= "010101";
                    when "0111010001010111" => rgb <= "010101";
                    when "0111010001011000" => rgb <= "010101";
                    when "0111010001011001" => rgb <= "010101";
                    when "0111010001011010" => rgb <= "010101";
                    when "0111010001011011" => rgb <= "010101";
                    when "0111010001011100" => rgb <= "010101";
                    when "0111010001011101" => rgb <= "010101";
                    when "0111010001011110" => rgb <= "010101";
                    when "0111010001100100" => rgb <= "010101";
                    when "0111010001100101" => rgb <= "010101";
                    when "0111010001100110" => rgb <= "010101";
                    when "0111010001100111" => rgb <= "010101";
                    when "0111010001101000" => rgb <= "010101";
                    when "0111010001101001" => rgb <= "010101";
                    when "0111010001101010" => rgb <= "010101";
                    when "0111010001101011" => rgb <= "010101";
                    when "0111010001101101" => rgb <= "010101";
                    when "0111010001101111" => rgb <= "010101";
                    when "0111010001110011" => rgb <= "010101";
                    when "0111010001110100" => rgb <= "010101";
                    when "0111010001110101" => rgb <= "010101";
                    when "0111010001110110" => rgb <= "010101";
                    when "0111010001110111" => rgb <= "010101";
                    when "0111010001111000" => rgb <= "010101";
                    when "0111010001111001" => rgb <= "010101";
                    when "0111010001111010" => rgb <= "010101";
                    when "0111010001111011" => rgb <= "010101";
                    when "0111010001111100" => rgb <= "010101";
                    when "0111010001111101" => rgb <= "010101";
                    when "0111010001111110" => rgb <= "010101";
                    when "0111010010000100" => rgb <= "010101";
                    when "0111010010001001" => rgb <= "010101";
                    when "0111010010001010" => rgb <= "010101";
                    when "0111010010001011" => rgb <= "010101";
                    when "0111010010001100" => rgb <= "010101";
                    when "0111010010001101" => rgb <= "010101";
                    when "0111010010001110" => rgb <= "010101";
                    when "0111010010010100" => rgb <= "010101";
                    when "0111010010011110" => rgb <= "010101";
                    when "0111010100000000" => rgb <= "101010";
                    when "0111010100000001" => rgb <= "101010";
                    when "0111010100000100" => rgb <= "010101";
                    when "0111010100000101" => rgb <= "010101";
                    when "0111010100000110" => rgb <= "010101";
                    when "0111010100000111" => rgb <= "010101";
                    when "0111010100001000" => rgb <= "010101";
                    when "0111010100001001" => rgb <= "010101";
                    when "0111010100001010" => rgb <= "010101";
                    when "0111010100001011" => rgb <= "010101";
                    when "0111010100001100" => rgb <= "010101";
                    when "0111010100010000" => rgb <= "101010";
                    when "0111010100010001" => rgb <= "101010";
                    when "0111010100010100" => rgb <= "010101";
                    when "0111010100010111" => rgb <= "010101";
                    when "0111010100011000" => rgb <= "010101";
                    when "0111010100011001" => rgb <= "010101";
                    when "0111010100011100" => rgb <= "010101";
                    when "0111010100100000" => rgb <= "101010";
                    when "0111010100100001" => rgb <= "101010";
                    when "0111010100100100" => rgb <= "010101";
                    when "0111010100101100" => rgb <= "010101";
                    when "0111010100110000" => rgb <= "101010";
                    when "0111010100110001" => rgb <= "101010";
                    when "0111010100110100" => rgb <= "010101";
                    when "0111010100110101" => rgb <= "010101";
                    when "0111010100110110" => rgb <= "010101";
                    when "0111010100110111" => rgb <= "010101";
                    when "0111010100111000" => rgb <= "010101";
                    when "0111010100111001" => rgb <= "010101";
                    when "0111010100111010" => rgb <= "010101";
                    when "0111010100111011" => rgb <= "010101";
                    when "0111010100111100" => rgb <= "010101";
                    when "0111010101000000" => rgb <= "101010";
                    when "0111010101000001" => rgb <= "101010";
                    when "0111010101000011" => rgb <= "010101";
                    when "0111010101000100" => rgb <= "010101";
                    when "0111010101000101" => rgb <= "010101";
                    when "0111010101000111" => rgb <= "010101";
                    when "0111010101001000" => rgb <= "010101";
                    when "0111010101001001" => rgb <= "010101";
                    when "0111010101001010" => rgb <= "010101";
                    when "0111010101001011" => rgb <= "010101";
                    when "0111010101001100" => rgb <= "010101";
                    when "0111010101001101" => rgb <= "010101";
                    when "0111010101010000" => rgb <= "101010";
                    when "0111010101010001" => rgb <= "101010";
                    when "0111010101010100" => rgb <= "010101";
                    when "0111010101010101" => rgb <= "010101";
                    when "0111010101010111" => rgb <= "010101";
                    when "0111010101011000" => rgb <= "101010";
                    when "0111010101011001" => rgb <= "010101";
                    when "0111010101011010" => rgb <= "010101";
                    when "0111010101011011" => rgb <= "010101";
                    when "0111010101011100" => rgb <= "010101";
                    when "0111010101011101" => rgb <= "010101";
                    when "0111010101100101" => rgb <= "010101";
                    when "0111010101100110" => rgb <= "010101";
                    when "0111010101100111" => rgb <= "010101";
                    when "0111010101101000" => rgb <= "010101";
                    when "0111010101101001" => rgb <= "010101";
                    when "0111010101101010" => rgb <= "010101";
                    when "0111010101101011" => rgb <= "010101";
                    when "0111010101101101" => rgb <= "010101";
                    when "0111010101101111" => rgb <= "010101";
                    when "0111010101110000" => rgb <= "101010";
                    when "0111010101110001" => rgb <= "101010";
                    when "0111010101110011" => rgb <= "010101";
                    when "0111010101110100" => rgb <= "010101";
                    when "0111010101110101" => rgb <= "010101";
                    when "0111010101110110" => rgb <= "010101";
                    when "0111010101110111" => rgb <= "010101";
                    when "0111010101111000" => rgb <= "010101";
                    when "0111010101111001" => rgb <= "010101";
                    when "0111010101111010" => rgb <= "010101";
                    when "0111010101111011" => rgb <= "010101";
                    when "0111010101111100" => rgb <= "010101";
                    when "0111010101111101" => rgb <= "010101";
                    when "0111010101111110" => rgb <= "010101";
                    when "0111010110000000" => rgb <= "101010";
                    when "0111010110000001" => rgb <= "101010";
                    when "0111010110000100" => rgb <= "010101";
                    when "0111010110001100" => rgb <= "010101";
                    when "0111010110001101" => rgb <= "010101";
                    when "0111010110001110" => rgb <= "010101";
                    when "0111010110010000" => rgb <= "101010";
                    when "0111010110010001" => rgb <= "101010";
                    when "0111010110010100" => rgb <= "010101";
                    when "0111010110011101" => rgb <= "010101";
                    when "0111010110011110" => rgb <= "010101";
                    when "0111011000000100" => rgb <= "010101";
                    when "0111011000000101" => rgb <= "010101";
                    when "0111011000000110" => rgb <= "010101";
                    when "0111011000000111" => rgb <= "010101";
                    when "0111011000001000" => rgb <= "010101";
                    when "0111011000001001" => rgb <= "010101";
                    when "0111011000001010" => rgb <= "010101";
                    when "0111011000001011" => rgb <= "010101";
                    when "0111011000001100" => rgb <= "010101";
                    when "0111011000001101" => rgb <= "010101";
                    when "0111011000010100" => rgb <= "010101";
                    when "0111011000010101" => rgb <= "010101";
                    when "0111011000010110" => rgb <= "010101";
                    when "0111011000010111" => rgb <= "010101";
                    when "0111011000011000" => rgb <= "010101";
                    when "0111011000011001" => rgb <= "010101";
                    when "0111011000011010" => rgb <= "010101";
                    when "0111011000011011" => rgb <= "010101";
                    when "0111011000011100" => rgb <= "010101";
                    when "0111011000011101" => rgb <= "010101";
                    when "0111011000100100" => rgb <= "010101";
                    when "0111011000100101" => rgb <= "010101";
                    when "0111011000100110" => rgb <= "010101";
                    when "0111011000100111" => rgb <= "010101";
                    when "0111011000101000" => rgb <= "010101";
                    when "0111011000101001" => rgb <= "010101";
                    when "0111011000101010" => rgb <= "010101";
                    when "0111011000101011" => rgb <= "010101";
                    when "0111011000101100" => rgb <= "010101";
                    when "0111011000101101" => rgb <= "010101";
                    when "0111011000110100" => rgb <= "010101";
                    when "0111011000110101" => rgb <= "010101";
                    when "0111011000110110" => rgb <= "010101";
                    when "0111011000110111" => rgb <= "010101";
                    when "0111011000111000" => rgb <= "010101";
                    when "0111011000111001" => rgb <= "010101";
                    when "0111011000111010" => rgb <= "010101";
                    when "0111011000111011" => rgb <= "010101";
                    when "0111011000111100" => rgb <= "010101";
                    when "0111011000111101" => rgb <= "010101";
                    when "0111011001000100" => rgb <= "010101";
                    when "0111011001000101" => rgb <= "010101";
                    when "0111011001000110" => rgb <= "010101";
                    when "0111011001000111" => rgb <= "010101";
                    when "0111011001001000" => rgb <= "010101";
                    when "0111011001001001" => rgb <= "010101";
                    when "0111011001001010" => rgb <= "010101";
                    when "0111011001001011" => rgb <= "010101";
                    when "0111011001001101" => rgb <= "010101";
                    when "0111011001010101" => rgb <= "010101";
                    when "0111011001010111" => rgb <= "010101";
                    when "0111011001011000" => rgb <= "101010";
                    when "0111011001011001" => rgb <= "010101";
                    when "0111011001011010" => rgb <= "010101";
                    when "0111011001011011" => rgb <= "010101";
                    when "0111011001011100" => rgb <= "010101";
                    when "0111011001011101" => rgb <= "010101";
                    when "0111011001100000" => rgb <= "010000";
                    when "0111011001100001" => rgb <= "010000";
                    when "0111011001100010" => rgb <= "010000";
                    when "0111011001100101" => rgb <= "010101";
                    when "0111011001100110" => rgb <= "010101";
                    when "0111011001100111" => rgb <= "010101";
                    when "0111011001101000" => rgb <= "010101";
                    when "0111011001101001" => rgb <= "010101";
                    when "0111011001101010" => rgb <= "010101";
                    when "0111011001101011" => rgb <= "010101";
                    when "0111011001101101" => rgb <= "010101";
                    when "0111011001101111" => rgb <= "010101";
                    when "0111011001110011" => rgb <= "010101";
                    when "0111011001110101" => rgb <= "010100";
                    when "0111011001110110" => rgb <= "010101";
                    when "0111011001110111" => rgb <= "010101";
                    when "0111011001111010" => rgb <= "010101";
                    when "0111011001111011" => rgb <= "010101";
                    when "0111011001111110" => rgb <= "010101";
                    when "0111011010000100" => rgb <= "010101";
                    when "0111011010000101" => rgb <= "010101";
                    when "0111011010000110" => rgb <= "010101";
                    when "0111011010000111" => rgb <= "010101";
                    when "0111011010001000" => rgb <= "010101";
                    when "0111011010001001" => rgb <= "010101";
                    when "0111011010001010" => rgb <= "010101";
                    when "0111011010001011" => rgb <= "010101";
                    when "0111011010001100" => rgb <= "010101";
                    when "0111011010001101" => rgb <= "010101";
                    when "0111011010001110" => rgb <= "010101";
                    when "0111011010010100" => rgb <= "010101";
                    when "0111011010010101" => rgb <= "010101";
                    when "0111011010010110" => rgb <= "010101";
                    when "0111011010010111" => rgb <= "010101";
                    when "0111011010011000" => rgb <= "010101";
                    when "0111011010011001" => rgb <= "010101";
                    when "0111011010011010" => rgb <= "010101";
                    when "0111011010011011" => rgb <= "010101";
                    when "0111011010011100" => rgb <= "010101";
                    when "0111011010011101" => rgb <= "010101";
                    when "0111011100000000" => rgb <= "101010";
                    when "0111011100000001" => rgb <= "101010";
                    when "0111011100010000" => rgb <= "101010";
                    when "0111011100010001" => rgb <= "101010";
                    when "0111011100100000" => rgb <= "101010";
                    when "0111011100100001" => rgb <= "101010";
                    when "0111011100110000" => rgb <= "101010";
                    when "0111011100110001" => rgb <= "101010";
                    when "0111011101000000" => rgb <= "101010";
                    when "0111011101000001" => rgb <= "101010";
                    when "0111011101010000" => rgb <= "101010";
                    when "0111011101010001" => rgb <= "101010";
                    when "0111011101010111" => rgb <= "010101";
                    when "0111011101011000" => rgb <= "101010";
                    when "0111011101011001" => rgb <= "010101";
                    when "0111011101011010" => rgb <= "010101";
                    when "0111011101011011" => rgb <= "010101";
                    when "0111011101011100" => rgb <= "010101";
                    when "0111011101011111" => rgb <= "010000";
                    when "0111011101100000" => rgb <= "010000";
                    when "0111011101100001" => rgb <= "010000";
                    when "0111011101100010" => rgb <= "010000";
                    when "0111011101100011" => rgb <= "010000";
                    when "0111011101100110" => rgb <= "010101";
                    when "0111011101100111" => rgb <= "010101";
                    when "0111011101101000" => rgb <= "010101";
                    when "0111011101101001" => rgb <= "010101";
                    when "0111011101101010" => rgb <= "010101";
                    when "0111011101101011" => rgb <= "010101";
                    when "0111011101110000" => rgb <= "101010";
                    when "0111011101110001" => rgb <= "101010";
                    when "0111011110000000" => rgb <= "101010";
                    when "0111011110000001" => rgb <= "101010";
                    when "0111011110010000" => rgb <= "101010";
                    when "0111011110010001" => rgb <= "101010";
                    when others => rgb <= "000000";
				end case;
			end if;
		end process;
end;